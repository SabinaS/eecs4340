`timescale 1ns/1ns
module spi_read (
	clk, rst
);

input clk, rst;

endmodule

