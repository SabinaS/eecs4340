`define display(A) $display("%s:%0d: %0d ns, cycle: %0d - %s", `__FILE__, `__LINE__, $time, $time / 20, $sformatf A );
