class transaction;
	/* ToDo */

endclass

class testing_env;

endclass

program ps2_tb (ps2_ifc.bench ds);

	transaction t;
	testing_env v;

endprogram
