`timescale 1ns/1ns
module sd_model_port (
          // spi_ifc.sdcard d
       );

// sdModel model (
// 				.spiClk(d.to_slave_o[0]),
// 				.spiDataIn(d.to_slave_o[1]),
// 				.spiDataOut(d.from_slave_i),
// 				.spiCS_n(d.to_slave_o[2])
// 			);

endmodule
