`timescale 1ns/1ns
module spi_read (
    to_slave_o, dat, valid_o, ready_o, ack_o,
    from_slave_i, read_i, write_i, valid_i, ready_i
);

endmodule

