`timescale 1ns/1ns

/* module for performing 4096 bit modular exponentiation */
module modexp(
	clk, rst, stall,
	exp, mod, key_i, start,
	key_o, done, valid
);
	input logic clk, rst, stall;
	input logic [4095:0] exp, mod; //would actually want to chunk this
	input logic [4095:0] key_i;
	input logic start;
	output logic [4095:0] key_o;
	output logic done, valid;


	logic [8191:0] intermediate;
	integer i;
	logic run;

	always_ff @(posedge clk) begin
		if(rst) begin
			run <= 1'b0;
			i <= 4095;
		end else if (!stall) begin
			if(start) begin
				run <= 1'b1;
			end
			if(run) begin
				if(i==0) begin
					i <= 4095;
					run <= 1'b0;
				end else begin
					i <= i-1;
				end
			end
		end
	end


	always_ff @(posedge clk) begin
		if(rst) begin
			intermediate <= 'b01;
			done <= 1'b0;
			valid <= 1'b0;
		end else if(!stall) begin
			if(run) begin
				if(i==0) begin
					key_o <= ((intermediate * (exp[i] ? key_i: 'b01)) % mod);
					done <= 1'b1;
					valid <= 1'b1;
				end else begin
					if (exp[i]) begin
						// intermediate <= (((intermediate * key_i) % mod) * ((intermediate * key_i) % mod)) % mod;
						intermediate <= (((intermediate * key_i) % mod) * ((intermediate * key_i) % mod)) % mod;
					end else begin
						intermediate <= (intermediate * intermediate) % mod;
					end
				end
			end
		end
	end

endmodule
