`timescale 1ns/1ns
// Multimedia File Encryption (Top Level)
module mfe (mfe_ifc.dut d);

    //TODO
    


    // // The PS/2 module wires (a small set for communication)
    // wire [15:0]         key_char_out;
    // wire                key_char_out_valid;
    
    // keyboard_driver keyboard (.char_o(key_char_out),
    //                         .char_valid_o(key_char_out_valid),
    //                         .clk(d.clk), .ps2_clk(d.ps2_clk),
    //                         .ps2_dat(d.ps2_dat));


endmodule
