`timescale 1ns/1ns

/* module for performing 4096 bit multiplication */
module multiplier2(
	clk, rst, a, b, o
);
	input logic clk, rst;
	input logic [4095:0] a, b; 
	output logic [4095:0] o;

	logic [8191:0] intermediate; 
	logic [11:0] stage; 

	assign o = intermediate[4095:0];


	always_ff @(posedge clk) begin
		if(rst) begin
			intermediate <= 'b0;
			stage <= 'b0;
		end else begin
			case(stage) 
12'd0: begin if(a[0]==1) 
	 		intermediate[4095+0:0+0] <= intermediate[4095+0:0+0] + a; end
12'd1: begin if(a[1]==1) 
	 		intermediate[4095+1:0+1] <= intermediate[4095+1:0+1] + a; end
12'd2: begin if(a[2]==1) 
	 		intermediate[4095+2:0+2] <= intermediate[4095+2:0+2] + a; end
12'd3: begin if(a[3]==1) 
	 		intermediate[4095+3:0+3] <= intermediate[4095+3:0+3] + a; end
12'd4: begin if(a[4]==1) 
	 		intermediate[4095+4:0+4] <= intermediate[4095+4:0+4] + a; end
12'd5: begin if(a[5]==1) 
	 		intermediate[4095+5:0+5] <= intermediate[4095+5:0+5] + a; end
12'd6: begin if(a[6]==1) 
	 		intermediate[4095+6:0+6] <= intermediate[4095+6:0+6] + a; end
12'd7: begin if(a[7]==1) 
	 		intermediate[4095+7:0+7] <= intermediate[4095+7:0+7] + a; end
12'd8: begin if(a[8]==1) 
	 		intermediate[4095+8:0+8] <= intermediate[4095+8:0+8] + a; end
12'd9: begin if(a[9]==1) 
	 		intermediate[4095+9:0+9] <= intermediate[4095+9:0+9] + a; end
12'd10: begin if(a[10]==1) 
	 		intermediate[4095+10:0+10] <= intermediate[4095+10:0+10] + a; end
12'd11: begin if(a[11]==1) 
	 		intermediate[4095+11:0+11] <= intermediate[4095+11:0+11] + a; end
12'd12: begin if(a[12]==1) 
	 		intermediate[4095+12:0+12] <= intermediate[4095+12:0+12] + a; end
12'd13: begin if(a[13]==1) 
	 		intermediate[4095+13:0+13] <= intermediate[4095+13:0+13] + a; end
12'd14: begin if(a[14]==1) 
	 		intermediate[4095+14:0+14] <= intermediate[4095+14:0+14] + a; end
12'd15: begin if(a[15]==1) 
	 		intermediate[4095+15:0+15] <= intermediate[4095+15:0+15] + a; end
12'd16: begin if(a[16]==1) 
	 		intermediate[4095+16:0+16] <= intermediate[4095+16:0+16] + a; end
12'd17: begin if(a[17]==1) 
	 		intermediate[4095+17:0+17] <= intermediate[4095+17:0+17] + a; end
12'd18: begin if(a[18]==1) 
	 		intermediate[4095+18:0+18] <= intermediate[4095+18:0+18] + a; end
12'd19: begin if(a[19]==1) 
	 		intermediate[4095+19:0+19] <= intermediate[4095+19:0+19] + a; end
12'd20: begin if(a[20]==1) 
	 		intermediate[4095+20:0+20] <= intermediate[4095+20:0+20] + a; end
12'd21: begin if(a[21]==1) 
	 		intermediate[4095+21:0+21] <= intermediate[4095+21:0+21] + a; end
12'd22: begin if(a[22]==1) 
	 		intermediate[4095+22:0+22] <= intermediate[4095+22:0+22] + a; end
12'd23: begin if(a[23]==1) 
	 		intermediate[4095+23:0+23] <= intermediate[4095+23:0+23] + a; end
12'd24: begin if(a[24]==1) 
	 		intermediate[4095+24:0+24] <= intermediate[4095+24:0+24] + a; end
12'd25: begin if(a[25]==1) 
	 		intermediate[4095+25:0+25] <= intermediate[4095+25:0+25] + a; end
12'd26: begin if(a[26]==1) 
	 		intermediate[4095+26:0+26] <= intermediate[4095+26:0+26] + a; end
12'd27: begin if(a[27]==1) 
	 		intermediate[4095+27:0+27] <= intermediate[4095+27:0+27] + a; end
12'd28: begin if(a[28]==1) 
	 		intermediate[4095+28:0+28] <= intermediate[4095+28:0+28] + a; end
12'd29: begin if(a[29]==1) 
	 		intermediate[4095+29:0+29] <= intermediate[4095+29:0+29] + a; end
12'd30: begin if(a[30]==1) 
	 		intermediate[4095+30:0+30] <= intermediate[4095+30:0+30] + a; end
12'd31: begin if(a[31]==1) 
	 		intermediate[4095+31:0+31] <= intermediate[4095+31:0+31] + a; end
12'd32: begin if(a[32]==1) 
	 		intermediate[4095+32:0+32] <= intermediate[4095+32:0+32] + a; end
12'd33: begin if(a[33]==1) 
	 		intermediate[4095+33:0+33] <= intermediate[4095+33:0+33] + a; end
12'd34: begin if(a[34]==1) 
	 		intermediate[4095+34:0+34] <= intermediate[4095+34:0+34] + a; end
12'd35: begin if(a[35]==1) 
	 		intermediate[4095+35:0+35] <= intermediate[4095+35:0+35] + a; end
12'd36: begin if(a[36]==1) 
	 		intermediate[4095+36:0+36] <= intermediate[4095+36:0+36] + a; end
12'd37: begin if(a[37]==1) 
	 		intermediate[4095+37:0+37] <= intermediate[4095+37:0+37] + a; end
12'd38: begin if(a[38]==1) 
	 		intermediate[4095+38:0+38] <= intermediate[4095+38:0+38] + a; end
12'd39: begin if(a[39]==1) 
	 		intermediate[4095+39:0+39] <= intermediate[4095+39:0+39] + a; end
12'd40: begin if(a[40]==1) 
	 		intermediate[4095+40:0+40] <= intermediate[4095+40:0+40] + a; end
12'd41: begin if(a[41]==1) 
	 		intermediate[4095+41:0+41] <= intermediate[4095+41:0+41] + a; end
12'd42: begin if(a[42]==1) 
	 		intermediate[4095+42:0+42] <= intermediate[4095+42:0+42] + a; end
12'd43: begin if(a[43]==1) 
	 		intermediate[4095+43:0+43] <= intermediate[4095+43:0+43] + a; end
12'd44: begin if(a[44]==1) 
	 		intermediate[4095+44:0+44] <= intermediate[4095+44:0+44] + a; end
12'd45: begin if(a[45]==1) 
	 		intermediate[4095+45:0+45] <= intermediate[4095+45:0+45] + a; end
12'd46: begin if(a[46]==1) 
	 		intermediate[4095+46:0+46] <= intermediate[4095+46:0+46] + a; end
12'd47: begin if(a[47]==1) 
	 		intermediate[4095+47:0+47] <= intermediate[4095+47:0+47] + a; end
12'd48: begin if(a[48]==1) 
	 		intermediate[4095+48:0+48] <= intermediate[4095+48:0+48] + a; end
12'd49: begin if(a[49]==1) 
	 		intermediate[4095+49:0+49] <= intermediate[4095+49:0+49] + a; end
12'd50: begin if(a[50]==1) 
	 		intermediate[4095+50:0+50] <= intermediate[4095+50:0+50] + a; end
12'd51: begin if(a[51]==1) 
	 		intermediate[4095+51:0+51] <= intermediate[4095+51:0+51] + a; end
12'd52: begin if(a[52]==1) 
	 		intermediate[4095+52:0+52] <= intermediate[4095+52:0+52] + a; end
12'd53: begin if(a[53]==1) 
	 		intermediate[4095+53:0+53] <= intermediate[4095+53:0+53] + a; end
12'd54: begin if(a[54]==1) 
	 		intermediate[4095+54:0+54] <= intermediate[4095+54:0+54] + a; end
12'd55: begin if(a[55]==1) 
	 		intermediate[4095+55:0+55] <= intermediate[4095+55:0+55] + a; end
12'd56: begin if(a[56]==1) 
	 		intermediate[4095+56:0+56] <= intermediate[4095+56:0+56] + a; end
12'd57: begin if(a[57]==1) 
	 		intermediate[4095+57:0+57] <= intermediate[4095+57:0+57] + a; end
12'd58: begin if(a[58]==1) 
	 		intermediate[4095+58:0+58] <= intermediate[4095+58:0+58] + a; end
12'd59: begin if(a[59]==1) 
	 		intermediate[4095+59:0+59] <= intermediate[4095+59:0+59] + a; end
12'd60: begin if(a[60]==1) 
	 		intermediate[4095+60:0+60] <= intermediate[4095+60:0+60] + a; end
12'd61: begin if(a[61]==1) 
	 		intermediate[4095+61:0+61] <= intermediate[4095+61:0+61] + a; end
12'd62: begin if(a[62]==1) 
	 		intermediate[4095+62:0+62] <= intermediate[4095+62:0+62] + a; end
12'd63: begin if(a[63]==1) 
	 		intermediate[4095+63:0+63] <= intermediate[4095+63:0+63] + a; end
12'd64: begin if(a[64]==1) 
	 		intermediate[4095+64:0+64] <= intermediate[4095+64:0+64] + a; end
12'd65: begin if(a[65]==1) 
	 		intermediate[4095+65:0+65] <= intermediate[4095+65:0+65] + a; end
12'd66: begin if(a[66]==1) 
	 		intermediate[4095+66:0+66] <= intermediate[4095+66:0+66] + a; end
12'd67: begin if(a[67]==1) 
	 		intermediate[4095+67:0+67] <= intermediate[4095+67:0+67] + a; end
12'd68: begin if(a[68]==1) 
	 		intermediate[4095+68:0+68] <= intermediate[4095+68:0+68] + a; end
12'd69: begin if(a[69]==1) 
	 		intermediate[4095+69:0+69] <= intermediate[4095+69:0+69] + a; end
12'd70: begin if(a[70]==1) 
	 		intermediate[4095+70:0+70] <= intermediate[4095+70:0+70] + a; end
12'd71: begin if(a[71]==1) 
	 		intermediate[4095+71:0+71] <= intermediate[4095+71:0+71] + a; end
12'd72: begin if(a[72]==1) 
	 		intermediate[4095+72:0+72] <= intermediate[4095+72:0+72] + a; end
12'd73: begin if(a[73]==1) 
	 		intermediate[4095+73:0+73] <= intermediate[4095+73:0+73] + a; end
12'd74: begin if(a[74]==1) 
	 		intermediate[4095+74:0+74] <= intermediate[4095+74:0+74] + a; end
12'd75: begin if(a[75]==1) 
	 		intermediate[4095+75:0+75] <= intermediate[4095+75:0+75] + a; end
12'd76: begin if(a[76]==1) 
	 		intermediate[4095+76:0+76] <= intermediate[4095+76:0+76] + a; end
12'd77: begin if(a[77]==1) 
	 		intermediate[4095+77:0+77] <= intermediate[4095+77:0+77] + a; end
12'd78: begin if(a[78]==1) 
	 		intermediate[4095+78:0+78] <= intermediate[4095+78:0+78] + a; end
12'd79: begin if(a[79]==1) 
	 		intermediate[4095+79:0+79] <= intermediate[4095+79:0+79] + a; end
12'd80: begin if(a[80]==1) 
	 		intermediate[4095+80:0+80] <= intermediate[4095+80:0+80] + a; end
12'd81: begin if(a[81]==1) 
	 		intermediate[4095+81:0+81] <= intermediate[4095+81:0+81] + a; end
12'd82: begin if(a[82]==1) 
	 		intermediate[4095+82:0+82] <= intermediate[4095+82:0+82] + a; end
12'd83: begin if(a[83]==1) 
	 		intermediate[4095+83:0+83] <= intermediate[4095+83:0+83] + a; end
12'd84: begin if(a[84]==1) 
	 		intermediate[4095+84:0+84] <= intermediate[4095+84:0+84] + a; end
12'd85: begin if(a[85]==1) 
	 		intermediate[4095+85:0+85] <= intermediate[4095+85:0+85] + a; end
12'd86: begin if(a[86]==1) 
	 		intermediate[4095+86:0+86] <= intermediate[4095+86:0+86] + a; end
12'd87: begin if(a[87]==1) 
	 		intermediate[4095+87:0+87] <= intermediate[4095+87:0+87] + a; end
12'd88: begin if(a[88]==1) 
	 		intermediate[4095+88:0+88] <= intermediate[4095+88:0+88] + a; end
12'd89: begin if(a[89]==1) 
	 		intermediate[4095+89:0+89] <= intermediate[4095+89:0+89] + a; end
12'd90: begin if(a[90]==1) 
	 		intermediate[4095+90:0+90] <= intermediate[4095+90:0+90] + a; end
12'd91: begin if(a[91]==1) 
	 		intermediate[4095+91:0+91] <= intermediate[4095+91:0+91] + a; end
12'd92: begin if(a[92]==1) 
	 		intermediate[4095+92:0+92] <= intermediate[4095+92:0+92] + a; end
12'd93: begin if(a[93]==1) 
	 		intermediate[4095+93:0+93] <= intermediate[4095+93:0+93] + a; end
12'd94: begin if(a[94]==1) 
	 		intermediate[4095+94:0+94] <= intermediate[4095+94:0+94] + a; end
12'd95: begin if(a[95]==1) 
	 		intermediate[4095+95:0+95] <= intermediate[4095+95:0+95] + a; end
12'd96: begin if(a[96]==1) 
	 		intermediate[4095+96:0+96] <= intermediate[4095+96:0+96] + a; end
12'd97: begin if(a[97]==1) 
	 		intermediate[4095+97:0+97] <= intermediate[4095+97:0+97] + a; end
12'd98: begin if(a[98]==1) 
	 		intermediate[4095+98:0+98] <= intermediate[4095+98:0+98] + a; end
12'd99: begin if(a[99]==1) 
	 		intermediate[4095+99:0+99] <= intermediate[4095+99:0+99] + a; end
12'd100: begin if(a[100]==1) 
	 		intermediate[4095+100:0+100] <= intermediate[4095+100:0+100] + a; end
12'd101: begin if(a[101]==1) 
	 		intermediate[4095+101:0+101] <= intermediate[4095+101:0+101] + a; end
12'd102: begin if(a[102]==1) 
	 		intermediate[4095+102:0+102] <= intermediate[4095+102:0+102] + a; end
12'd103: begin if(a[103]==1) 
	 		intermediate[4095+103:0+103] <= intermediate[4095+103:0+103] + a; end
12'd104: begin if(a[104]==1) 
	 		intermediate[4095+104:0+104] <= intermediate[4095+104:0+104] + a; end
12'd105: begin if(a[105]==1) 
	 		intermediate[4095+105:0+105] <= intermediate[4095+105:0+105] + a; end
12'd106: begin if(a[106]==1) 
	 		intermediate[4095+106:0+106] <= intermediate[4095+106:0+106] + a; end
12'd107: begin if(a[107]==1) 
	 		intermediate[4095+107:0+107] <= intermediate[4095+107:0+107] + a; end
12'd108: begin if(a[108]==1) 
	 		intermediate[4095+108:0+108] <= intermediate[4095+108:0+108] + a; end
12'd109: begin if(a[109]==1) 
	 		intermediate[4095+109:0+109] <= intermediate[4095+109:0+109] + a; end
12'd110: begin if(a[110]==1) 
	 		intermediate[4095+110:0+110] <= intermediate[4095+110:0+110] + a; end
12'd111: begin if(a[111]==1) 
	 		intermediate[4095+111:0+111] <= intermediate[4095+111:0+111] + a; end
12'd112: begin if(a[112]==1) 
	 		intermediate[4095+112:0+112] <= intermediate[4095+112:0+112] + a; end
12'd113: begin if(a[113]==1) 
	 		intermediate[4095+113:0+113] <= intermediate[4095+113:0+113] + a; end
12'd114: begin if(a[114]==1) 
	 		intermediate[4095+114:0+114] <= intermediate[4095+114:0+114] + a; end
12'd115: begin if(a[115]==1) 
	 		intermediate[4095+115:0+115] <= intermediate[4095+115:0+115] + a; end
12'd116: begin if(a[116]==1) 
	 		intermediate[4095+116:0+116] <= intermediate[4095+116:0+116] + a; end
12'd117: begin if(a[117]==1) 
	 		intermediate[4095+117:0+117] <= intermediate[4095+117:0+117] + a; end
12'd118: begin if(a[118]==1) 
	 		intermediate[4095+118:0+118] <= intermediate[4095+118:0+118] + a; end
12'd119: begin if(a[119]==1) 
	 		intermediate[4095+119:0+119] <= intermediate[4095+119:0+119] + a; end
12'd120: begin if(a[120]==1) 
	 		intermediate[4095+120:0+120] <= intermediate[4095+120:0+120] + a; end
12'd121: begin if(a[121]==1) 
	 		intermediate[4095+121:0+121] <= intermediate[4095+121:0+121] + a; end
12'd122: begin if(a[122]==1) 
	 		intermediate[4095+122:0+122] <= intermediate[4095+122:0+122] + a; end
12'd123: begin if(a[123]==1) 
	 		intermediate[4095+123:0+123] <= intermediate[4095+123:0+123] + a; end
12'd124: begin if(a[124]==1) 
	 		intermediate[4095+124:0+124] <= intermediate[4095+124:0+124] + a; end
12'd125: begin if(a[125]==1) 
	 		intermediate[4095+125:0+125] <= intermediate[4095+125:0+125] + a; end
12'd126: begin if(a[126]==1) 
	 		intermediate[4095+126:0+126] <= intermediate[4095+126:0+126] + a; end
12'd127: begin if(a[127]==1) 
	 		intermediate[4095+127:0+127] <= intermediate[4095+127:0+127] + a; end
12'd128: begin if(a[128]==1) 
	 		intermediate[4095+128:0+128] <= intermediate[4095+128:0+128] + a; end
12'd129: begin if(a[129]==1) 
	 		intermediate[4095+129:0+129] <= intermediate[4095+129:0+129] + a; end
12'd130: begin if(a[130]==1) 
	 		intermediate[4095+130:0+130] <= intermediate[4095+130:0+130] + a; end
12'd131: begin if(a[131]==1) 
	 		intermediate[4095+131:0+131] <= intermediate[4095+131:0+131] + a; end
12'd132: begin if(a[132]==1) 
	 		intermediate[4095+132:0+132] <= intermediate[4095+132:0+132] + a; end
12'd133: begin if(a[133]==1) 
	 		intermediate[4095+133:0+133] <= intermediate[4095+133:0+133] + a; end
12'd134: begin if(a[134]==1) 
	 		intermediate[4095+134:0+134] <= intermediate[4095+134:0+134] + a; end
12'd135: begin if(a[135]==1) 
	 		intermediate[4095+135:0+135] <= intermediate[4095+135:0+135] + a; end
12'd136: begin if(a[136]==1) 
	 		intermediate[4095+136:0+136] <= intermediate[4095+136:0+136] + a; end
12'd137: begin if(a[137]==1) 
	 		intermediate[4095+137:0+137] <= intermediate[4095+137:0+137] + a; end
12'd138: begin if(a[138]==1) 
	 		intermediate[4095+138:0+138] <= intermediate[4095+138:0+138] + a; end
12'd139: begin if(a[139]==1) 
	 		intermediate[4095+139:0+139] <= intermediate[4095+139:0+139] + a; end
12'd140: begin if(a[140]==1) 
	 		intermediate[4095+140:0+140] <= intermediate[4095+140:0+140] + a; end
12'd141: begin if(a[141]==1) 
	 		intermediate[4095+141:0+141] <= intermediate[4095+141:0+141] + a; end
12'd142: begin if(a[142]==1) 
	 		intermediate[4095+142:0+142] <= intermediate[4095+142:0+142] + a; end
12'd143: begin if(a[143]==1) 
	 		intermediate[4095+143:0+143] <= intermediate[4095+143:0+143] + a; end
12'd144: begin if(a[144]==1) 
	 		intermediate[4095+144:0+144] <= intermediate[4095+144:0+144] + a; end
12'd145: begin if(a[145]==1) 
	 		intermediate[4095+145:0+145] <= intermediate[4095+145:0+145] + a; end
12'd146: begin if(a[146]==1) 
	 		intermediate[4095+146:0+146] <= intermediate[4095+146:0+146] + a; end
12'd147: begin if(a[147]==1) 
	 		intermediate[4095+147:0+147] <= intermediate[4095+147:0+147] + a; end
12'd148: begin if(a[148]==1) 
	 		intermediate[4095+148:0+148] <= intermediate[4095+148:0+148] + a; end
12'd149: begin if(a[149]==1) 
	 		intermediate[4095+149:0+149] <= intermediate[4095+149:0+149] + a; end
12'd150: begin if(a[150]==1) 
	 		intermediate[4095+150:0+150] <= intermediate[4095+150:0+150] + a; end
12'd151: begin if(a[151]==1) 
	 		intermediate[4095+151:0+151] <= intermediate[4095+151:0+151] + a; end
12'd152: begin if(a[152]==1) 
	 		intermediate[4095+152:0+152] <= intermediate[4095+152:0+152] + a; end
12'd153: begin if(a[153]==1) 
	 		intermediate[4095+153:0+153] <= intermediate[4095+153:0+153] + a; end
12'd154: begin if(a[154]==1) 
	 		intermediate[4095+154:0+154] <= intermediate[4095+154:0+154] + a; end
12'd155: begin if(a[155]==1) 
	 		intermediate[4095+155:0+155] <= intermediate[4095+155:0+155] + a; end
12'd156: begin if(a[156]==1) 
	 		intermediate[4095+156:0+156] <= intermediate[4095+156:0+156] + a; end
12'd157: begin if(a[157]==1) 
	 		intermediate[4095+157:0+157] <= intermediate[4095+157:0+157] + a; end
12'd158: begin if(a[158]==1) 
	 		intermediate[4095+158:0+158] <= intermediate[4095+158:0+158] + a; end
12'd159: begin if(a[159]==1) 
	 		intermediate[4095+159:0+159] <= intermediate[4095+159:0+159] + a; end
12'd160: begin if(a[160]==1) 
	 		intermediate[4095+160:0+160] <= intermediate[4095+160:0+160] + a; end
12'd161: begin if(a[161]==1) 
	 		intermediate[4095+161:0+161] <= intermediate[4095+161:0+161] + a; end
12'd162: begin if(a[162]==1) 
	 		intermediate[4095+162:0+162] <= intermediate[4095+162:0+162] + a; end
12'd163: begin if(a[163]==1) 
	 		intermediate[4095+163:0+163] <= intermediate[4095+163:0+163] + a; end
12'd164: begin if(a[164]==1) 
	 		intermediate[4095+164:0+164] <= intermediate[4095+164:0+164] + a; end
12'd165: begin if(a[165]==1) 
	 		intermediate[4095+165:0+165] <= intermediate[4095+165:0+165] + a; end
12'd166: begin if(a[166]==1) 
	 		intermediate[4095+166:0+166] <= intermediate[4095+166:0+166] + a; end
12'd167: begin if(a[167]==1) 
	 		intermediate[4095+167:0+167] <= intermediate[4095+167:0+167] + a; end
12'd168: begin if(a[168]==1) 
	 		intermediate[4095+168:0+168] <= intermediate[4095+168:0+168] + a; end
12'd169: begin if(a[169]==1) 
	 		intermediate[4095+169:0+169] <= intermediate[4095+169:0+169] + a; end
12'd170: begin if(a[170]==1) 
	 		intermediate[4095+170:0+170] <= intermediate[4095+170:0+170] + a; end
12'd171: begin if(a[171]==1) 
	 		intermediate[4095+171:0+171] <= intermediate[4095+171:0+171] + a; end
12'd172: begin if(a[172]==1) 
	 		intermediate[4095+172:0+172] <= intermediate[4095+172:0+172] + a; end
12'd173: begin if(a[173]==1) 
	 		intermediate[4095+173:0+173] <= intermediate[4095+173:0+173] + a; end
12'd174: begin if(a[174]==1) 
	 		intermediate[4095+174:0+174] <= intermediate[4095+174:0+174] + a; end
12'd175: begin if(a[175]==1) 
	 		intermediate[4095+175:0+175] <= intermediate[4095+175:0+175] + a; end
12'd176: begin if(a[176]==1) 
	 		intermediate[4095+176:0+176] <= intermediate[4095+176:0+176] + a; end
12'd177: begin if(a[177]==1) 
	 		intermediate[4095+177:0+177] <= intermediate[4095+177:0+177] + a; end
12'd178: begin if(a[178]==1) 
	 		intermediate[4095+178:0+178] <= intermediate[4095+178:0+178] + a; end
12'd179: begin if(a[179]==1) 
	 		intermediate[4095+179:0+179] <= intermediate[4095+179:0+179] + a; end
12'd180: begin if(a[180]==1) 
	 		intermediate[4095+180:0+180] <= intermediate[4095+180:0+180] + a; end
12'd181: begin if(a[181]==1) 
	 		intermediate[4095+181:0+181] <= intermediate[4095+181:0+181] + a; end
12'd182: begin if(a[182]==1) 
	 		intermediate[4095+182:0+182] <= intermediate[4095+182:0+182] + a; end
12'd183: begin if(a[183]==1) 
	 		intermediate[4095+183:0+183] <= intermediate[4095+183:0+183] + a; end
12'd184: begin if(a[184]==1) 
	 		intermediate[4095+184:0+184] <= intermediate[4095+184:0+184] + a; end
12'd185: begin if(a[185]==1) 
	 		intermediate[4095+185:0+185] <= intermediate[4095+185:0+185] + a; end
12'd186: begin if(a[186]==1) 
	 		intermediate[4095+186:0+186] <= intermediate[4095+186:0+186] + a; end
12'd187: begin if(a[187]==1) 
	 		intermediate[4095+187:0+187] <= intermediate[4095+187:0+187] + a; end
12'd188: begin if(a[188]==1) 
	 		intermediate[4095+188:0+188] <= intermediate[4095+188:0+188] + a; end
12'd189: begin if(a[189]==1) 
	 		intermediate[4095+189:0+189] <= intermediate[4095+189:0+189] + a; end
12'd190: begin if(a[190]==1) 
	 		intermediate[4095+190:0+190] <= intermediate[4095+190:0+190] + a; end
12'd191: begin if(a[191]==1) 
	 		intermediate[4095+191:0+191] <= intermediate[4095+191:0+191] + a; end
12'd192: begin if(a[192]==1) 
	 		intermediate[4095+192:0+192] <= intermediate[4095+192:0+192] + a; end
12'd193: begin if(a[193]==1) 
	 		intermediate[4095+193:0+193] <= intermediate[4095+193:0+193] + a; end
12'd194: begin if(a[194]==1) 
	 		intermediate[4095+194:0+194] <= intermediate[4095+194:0+194] + a; end
12'd195: begin if(a[195]==1) 
	 		intermediate[4095+195:0+195] <= intermediate[4095+195:0+195] + a; end
12'd196: begin if(a[196]==1) 
	 		intermediate[4095+196:0+196] <= intermediate[4095+196:0+196] + a; end
12'd197: begin if(a[197]==1) 
	 		intermediate[4095+197:0+197] <= intermediate[4095+197:0+197] + a; end
12'd198: begin if(a[198]==1) 
	 		intermediate[4095+198:0+198] <= intermediate[4095+198:0+198] + a; end
12'd199: begin if(a[199]==1) 
	 		intermediate[4095+199:0+199] <= intermediate[4095+199:0+199] + a; end
12'd200: begin if(a[200]==1) 
	 		intermediate[4095+200:0+200] <= intermediate[4095+200:0+200] + a; end
12'd201: begin if(a[201]==1) 
	 		intermediate[4095+201:0+201] <= intermediate[4095+201:0+201] + a; end
12'd202: begin if(a[202]==1) 
	 		intermediate[4095+202:0+202] <= intermediate[4095+202:0+202] + a; end
12'd203: begin if(a[203]==1) 
	 		intermediate[4095+203:0+203] <= intermediate[4095+203:0+203] + a; end
12'd204: begin if(a[204]==1) 
	 		intermediate[4095+204:0+204] <= intermediate[4095+204:0+204] + a; end
12'd205: begin if(a[205]==1) 
	 		intermediate[4095+205:0+205] <= intermediate[4095+205:0+205] + a; end
12'd206: begin if(a[206]==1) 
	 		intermediate[4095+206:0+206] <= intermediate[4095+206:0+206] + a; end
12'd207: begin if(a[207]==1) 
	 		intermediate[4095+207:0+207] <= intermediate[4095+207:0+207] + a; end
12'd208: begin if(a[208]==1) 
	 		intermediate[4095+208:0+208] <= intermediate[4095+208:0+208] + a; end
12'd209: begin if(a[209]==1) 
	 		intermediate[4095+209:0+209] <= intermediate[4095+209:0+209] + a; end
12'd210: begin if(a[210]==1) 
	 		intermediate[4095+210:0+210] <= intermediate[4095+210:0+210] + a; end
12'd211: begin if(a[211]==1) 
	 		intermediate[4095+211:0+211] <= intermediate[4095+211:0+211] + a; end
12'd212: begin if(a[212]==1) 
	 		intermediate[4095+212:0+212] <= intermediate[4095+212:0+212] + a; end
12'd213: begin if(a[213]==1) 
	 		intermediate[4095+213:0+213] <= intermediate[4095+213:0+213] + a; end
12'd214: begin if(a[214]==1) 
	 		intermediate[4095+214:0+214] <= intermediate[4095+214:0+214] + a; end
12'd215: begin if(a[215]==1) 
	 		intermediate[4095+215:0+215] <= intermediate[4095+215:0+215] + a; end
12'd216: begin if(a[216]==1) 
	 		intermediate[4095+216:0+216] <= intermediate[4095+216:0+216] + a; end
12'd217: begin if(a[217]==1) 
	 		intermediate[4095+217:0+217] <= intermediate[4095+217:0+217] + a; end
12'd218: begin if(a[218]==1) 
	 		intermediate[4095+218:0+218] <= intermediate[4095+218:0+218] + a; end
12'd219: begin if(a[219]==1) 
	 		intermediate[4095+219:0+219] <= intermediate[4095+219:0+219] + a; end
12'd220: begin if(a[220]==1) 
	 		intermediate[4095+220:0+220] <= intermediate[4095+220:0+220] + a; end
12'd221: begin if(a[221]==1) 
	 		intermediate[4095+221:0+221] <= intermediate[4095+221:0+221] + a; end
12'd222: begin if(a[222]==1) 
	 		intermediate[4095+222:0+222] <= intermediate[4095+222:0+222] + a; end
12'd223: begin if(a[223]==1) 
	 		intermediate[4095+223:0+223] <= intermediate[4095+223:0+223] + a; end
12'd224: begin if(a[224]==1) 
	 		intermediate[4095+224:0+224] <= intermediate[4095+224:0+224] + a; end
12'd225: begin if(a[225]==1) 
	 		intermediate[4095+225:0+225] <= intermediate[4095+225:0+225] + a; end
12'd226: begin if(a[226]==1) 
	 		intermediate[4095+226:0+226] <= intermediate[4095+226:0+226] + a; end
12'd227: begin if(a[227]==1) 
	 		intermediate[4095+227:0+227] <= intermediate[4095+227:0+227] + a; end
12'd228: begin if(a[228]==1) 
	 		intermediate[4095+228:0+228] <= intermediate[4095+228:0+228] + a; end
12'd229: begin if(a[229]==1) 
	 		intermediate[4095+229:0+229] <= intermediate[4095+229:0+229] + a; end
12'd230: begin if(a[230]==1) 
	 		intermediate[4095+230:0+230] <= intermediate[4095+230:0+230] + a; end
12'd231: begin if(a[231]==1) 
	 		intermediate[4095+231:0+231] <= intermediate[4095+231:0+231] + a; end
12'd232: begin if(a[232]==1) 
	 		intermediate[4095+232:0+232] <= intermediate[4095+232:0+232] + a; end
12'd233: begin if(a[233]==1) 
	 		intermediate[4095+233:0+233] <= intermediate[4095+233:0+233] + a; end
12'd234: begin if(a[234]==1) 
	 		intermediate[4095+234:0+234] <= intermediate[4095+234:0+234] + a; end
12'd235: begin if(a[235]==1) 
	 		intermediate[4095+235:0+235] <= intermediate[4095+235:0+235] + a; end
12'd236: begin if(a[236]==1) 
	 		intermediate[4095+236:0+236] <= intermediate[4095+236:0+236] + a; end
12'd237: begin if(a[237]==1) 
	 		intermediate[4095+237:0+237] <= intermediate[4095+237:0+237] + a; end
12'd238: begin if(a[238]==1) 
	 		intermediate[4095+238:0+238] <= intermediate[4095+238:0+238] + a; end
12'd239: begin if(a[239]==1) 
	 		intermediate[4095+239:0+239] <= intermediate[4095+239:0+239] + a; end
12'd240: begin if(a[240]==1) 
	 		intermediate[4095+240:0+240] <= intermediate[4095+240:0+240] + a; end
12'd241: begin if(a[241]==1) 
	 		intermediate[4095+241:0+241] <= intermediate[4095+241:0+241] + a; end
12'd242: begin if(a[242]==1) 
	 		intermediate[4095+242:0+242] <= intermediate[4095+242:0+242] + a; end
12'd243: begin if(a[243]==1) 
	 		intermediate[4095+243:0+243] <= intermediate[4095+243:0+243] + a; end
12'd244: begin if(a[244]==1) 
	 		intermediate[4095+244:0+244] <= intermediate[4095+244:0+244] + a; end
12'd245: begin if(a[245]==1) 
	 		intermediate[4095+245:0+245] <= intermediate[4095+245:0+245] + a; end
12'd246: begin if(a[246]==1) 
	 		intermediate[4095+246:0+246] <= intermediate[4095+246:0+246] + a; end
12'd247: begin if(a[247]==1) 
	 		intermediate[4095+247:0+247] <= intermediate[4095+247:0+247] + a; end
12'd248: begin if(a[248]==1) 
	 		intermediate[4095+248:0+248] <= intermediate[4095+248:0+248] + a; end
12'd249: begin if(a[249]==1) 
	 		intermediate[4095+249:0+249] <= intermediate[4095+249:0+249] + a; end
12'd250: begin if(a[250]==1) 
	 		intermediate[4095+250:0+250] <= intermediate[4095+250:0+250] + a; end
12'd251: begin if(a[251]==1) 
	 		intermediate[4095+251:0+251] <= intermediate[4095+251:0+251] + a; end
12'd252: begin if(a[252]==1) 
	 		intermediate[4095+252:0+252] <= intermediate[4095+252:0+252] + a; end
12'd253: begin if(a[253]==1) 
	 		intermediate[4095+253:0+253] <= intermediate[4095+253:0+253] + a; end
12'd254: begin if(a[254]==1) 
	 		intermediate[4095+254:0+254] <= intermediate[4095+254:0+254] + a; end
12'd255: begin if(a[255]==1) 
	 		intermediate[4095+255:0+255] <= intermediate[4095+255:0+255] + a; end
12'd256: begin if(a[256]==1) 
	 		intermediate[4095+256:0+256] <= intermediate[4095+256:0+256] + a; end
12'd257: begin if(a[257]==1) 
	 		intermediate[4095+257:0+257] <= intermediate[4095+257:0+257] + a; end
12'd258: begin if(a[258]==1) 
	 		intermediate[4095+258:0+258] <= intermediate[4095+258:0+258] + a; end
12'd259: begin if(a[259]==1) 
	 		intermediate[4095+259:0+259] <= intermediate[4095+259:0+259] + a; end
12'd260: begin if(a[260]==1) 
	 		intermediate[4095+260:0+260] <= intermediate[4095+260:0+260] + a; end
12'd261: begin if(a[261]==1) 
	 		intermediate[4095+261:0+261] <= intermediate[4095+261:0+261] + a; end
12'd262: begin if(a[262]==1) 
	 		intermediate[4095+262:0+262] <= intermediate[4095+262:0+262] + a; end
12'd263: begin if(a[263]==1) 
	 		intermediate[4095+263:0+263] <= intermediate[4095+263:0+263] + a; end
12'd264: begin if(a[264]==1) 
	 		intermediate[4095+264:0+264] <= intermediate[4095+264:0+264] + a; end
12'd265: begin if(a[265]==1) 
	 		intermediate[4095+265:0+265] <= intermediate[4095+265:0+265] + a; end
12'd266: begin if(a[266]==1) 
	 		intermediate[4095+266:0+266] <= intermediate[4095+266:0+266] + a; end
12'd267: begin if(a[267]==1) 
	 		intermediate[4095+267:0+267] <= intermediate[4095+267:0+267] + a; end
12'd268: begin if(a[268]==1) 
	 		intermediate[4095+268:0+268] <= intermediate[4095+268:0+268] + a; end
12'd269: begin if(a[269]==1) 
	 		intermediate[4095+269:0+269] <= intermediate[4095+269:0+269] + a; end
12'd270: begin if(a[270]==1) 
	 		intermediate[4095+270:0+270] <= intermediate[4095+270:0+270] + a; end
12'd271: begin if(a[271]==1) 
	 		intermediate[4095+271:0+271] <= intermediate[4095+271:0+271] + a; end
12'd272: begin if(a[272]==1) 
	 		intermediate[4095+272:0+272] <= intermediate[4095+272:0+272] + a; end
12'd273: begin if(a[273]==1) 
	 		intermediate[4095+273:0+273] <= intermediate[4095+273:0+273] + a; end
12'd274: begin if(a[274]==1) 
	 		intermediate[4095+274:0+274] <= intermediate[4095+274:0+274] + a; end
12'd275: begin if(a[275]==1) 
	 		intermediate[4095+275:0+275] <= intermediate[4095+275:0+275] + a; end
12'd276: begin if(a[276]==1) 
	 		intermediate[4095+276:0+276] <= intermediate[4095+276:0+276] + a; end
12'd277: begin if(a[277]==1) 
	 		intermediate[4095+277:0+277] <= intermediate[4095+277:0+277] + a; end
12'd278: begin if(a[278]==1) 
	 		intermediate[4095+278:0+278] <= intermediate[4095+278:0+278] + a; end
12'd279: begin if(a[279]==1) 
	 		intermediate[4095+279:0+279] <= intermediate[4095+279:0+279] + a; end
12'd280: begin if(a[280]==1) 
	 		intermediate[4095+280:0+280] <= intermediate[4095+280:0+280] + a; end
12'd281: begin if(a[281]==1) 
	 		intermediate[4095+281:0+281] <= intermediate[4095+281:0+281] + a; end
12'd282: begin if(a[282]==1) 
	 		intermediate[4095+282:0+282] <= intermediate[4095+282:0+282] + a; end
12'd283: begin if(a[283]==1) 
	 		intermediate[4095+283:0+283] <= intermediate[4095+283:0+283] + a; end
12'd284: begin if(a[284]==1) 
	 		intermediate[4095+284:0+284] <= intermediate[4095+284:0+284] + a; end
12'd285: begin if(a[285]==1) 
	 		intermediate[4095+285:0+285] <= intermediate[4095+285:0+285] + a; end
12'd286: begin if(a[286]==1) 
	 		intermediate[4095+286:0+286] <= intermediate[4095+286:0+286] + a; end
12'd287: begin if(a[287]==1) 
	 		intermediate[4095+287:0+287] <= intermediate[4095+287:0+287] + a; end
12'd288: begin if(a[288]==1) 
	 		intermediate[4095+288:0+288] <= intermediate[4095+288:0+288] + a; end
12'd289: begin if(a[289]==1) 
	 		intermediate[4095+289:0+289] <= intermediate[4095+289:0+289] + a; end
12'd290: begin if(a[290]==1) 
	 		intermediate[4095+290:0+290] <= intermediate[4095+290:0+290] + a; end
12'd291: begin if(a[291]==1) 
	 		intermediate[4095+291:0+291] <= intermediate[4095+291:0+291] + a; end
12'd292: begin if(a[292]==1) 
	 		intermediate[4095+292:0+292] <= intermediate[4095+292:0+292] + a; end
12'd293: begin if(a[293]==1) 
	 		intermediate[4095+293:0+293] <= intermediate[4095+293:0+293] + a; end
12'd294: begin if(a[294]==1) 
	 		intermediate[4095+294:0+294] <= intermediate[4095+294:0+294] + a; end
12'd295: begin if(a[295]==1) 
	 		intermediate[4095+295:0+295] <= intermediate[4095+295:0+295] + a; end
12'd296: begin if(a[296]==1) 
	 		intermediate[4095+296:0+296] <= intermediate[4095+296:0+296] + a; end
12'd297: begin if(a[297]==1) 
	 		intermediate[4095+297:0+297] <= intermediate[4095+297:0+297] + a; end
12'd298: begin if(a[298]==1) 
	 		intermediate[4095+298:0+298] <= intermediate[4095+298:0+298] + a; end
12'd299: begin if(a[299]==1) 
	 		intermediate[4095+299:0+299] <= intermediate[4095+299:0+299] + a; end
12'd300: begin if(a[300]==1) 
	 		intermediate[4095+300:0+300] <= intermediate[4095+300:0+300] + a; end
12'd301: begin if(a[301]==1) 
	 		intermediate[4095+301:0+301] <= intermediate[4095+301:0+301] + a; end
12'd302: begin if(a[302]==1) 
	 		intermediate[4095+302:0+302] <= intermediate[4095+302:0+302] + a; end
12'd303: begin if(a[303]==1) 
	 		intermediate[4095+303:0+303] <= intermediate[4095+303:0+303] + a; end
12'd304: begin if(a[304]==1) 
	 		intermediate[4095+304:0+304] <= intermediate[4095+304:0+304] + a; end
12'd305: begin if(a[305]==1) 
	 		intermediate[4095+305:0+305] <= intermediate[4095+305:0+305] + a; end
12'd306: begin if(a[306]==1) 
	 		intermediate[4095+306:0+306] <= intermediate[4095+306:0+306] + a; end
12'd307: begin if(a[307]==1) 
	 		intermediate[4095+307:0+307] <= intermediate[4095+307:0+307] + a; end
12'd308: begin if(a[308]==1) 
	 		intermediate[4095+308:0+308] <= intermediate[4095+308:0+308] + a; end
12'd309: begin if(a[309]==1) 
	 		intermediate[4095+309:0+309] <= intermediate[4095+309:0+309] + a; end
12'd310: begin if(a[310]==1) 
	 		intermediate[4095+310:0+310] <= intermediate[4095+310:0+310] + a; end
12'd311: begin if(a[311]==1) 
	 		intermediate[4095+311:0+311] <= intermediate[4095+311:0+311] + a; end
12'd312: begin if(a[312]==1) 
	 		intermediate[4095+312:0+312] <= intermediate[4095+312:0+312] + a; end
12'd313: begin if(a[313]==1) 
	 		intermediate[4095+313:0+313] <= intermediate[4095+313:0+313] + a; end
12'd314: begin if(a[314]==1) 
	 		intermediate[4095+314:0+314] <= intermediate[4095+314:0+314] + a; end
12'd315: begin if(a[315]==1) 
	 		intermediate[4095+315:0+315] <= intermediate[4095+315:0+315] + a; end
12'd316: begin if(a[316]==1) 
	 		intermediate[4095+316:0+316] <= intermediate[4095+316:0+316] + a; end
12'd317: begin if(a[317]==1) 
	 		intermediate[4095+317:0+317] <= intermediate[4095+317:0+317] + a; end
12'd318: begin if(a[318]==1) 
	 		intermediate[4095+318:0+318] <= intermediate[4095+318:0+318] + a; end
12'd319: begin if(a[319]==1) 
	 		intermediate[4095+319:0+319] <= intermediate[4095+319:0+319] + a; end
12'd320: begin if(a[320]==1) 
	 		intermediate[4095+320:0+320] <= intermediate[4095+320:0+320] + a; end
12'd321: begin if(a[321]==1) 
	 		intermediate[4095+321:0+321] <= intermediate[4095+321:0+321] + a; end
12'd322: begin if(a[322]==1) 
	 		intermediate[4095+322:0+322] <= intermediate[4095+322:0+322] + a; end
12'd323: begin if(a[323]==1) 
	 		intermediate[4095+323:0+323] <= intermediate[4095+323:0+323] + a; end
12'd324: begin if(a[324]==1) 
	 		intermediate[4095+324:0+324] <= intermediate[4095+324:0+324] + a; end
12'd325: begin if(a[325]==1) 
	 		intermediate[4095+325:0+325] <= intermediate[4095+325:0+325] + a; end
12'd326: begin if(a[326]==1) 
	 		intermediate[4095+326:0+326] <= intermediate[4095+326:0+326] + a; end
12'd327: begin if(a[327]==1) 
	 		intermediate[4095+327:0+327] <= intermediate[4095+327:0+327] + a; end
12'd328: begin if(a[328]==1) 
	 		intermediate[4095+328:0+328] <= intermediate[4095+328:0+328] + a; end
12'd329: begin if(a[329]==1) 
	 		intermediate[4095+329:0+329] <= intermediate[4095+329:0+329] + a; end
12'd330: begin if(a[330]==1) 
	 		intermediate[4095+330:0+330] <= intermediate[4095+330:0+330] + a; end
12'd331: begin if(a[331]==1) 
	 		intermediate[4095+331:0+331] <= intermediate[4095+331:0+331] + a; end
12'd332: begin if(a[332]==1) 
	 		intermediate[4095+332:0+332] <= intermediate[4095+332:0+332] + a; end
12'd333: begin if(a[333]==1) 
	 		intermediate[4095+333:0+333] <= intermediate[4095+333:0+333] + a; end
12'd334: begin if(a[334]==1) 
	 		intermediate[4095+334:0+334] <= intermediate[4095+334:0+334] + a; end
12'd335: begin if(a[335]==1) 
	 		intermediate[4095+335:0+335] <= intermediate[4095+335:0+335] + a; end
12'd336: begin if(a[336]==1) 
	 		intermediate[4095+336:0+336] <= intermediate[4095+336:0+336] + a; end
12'd337: begin if(a[337]==1) 
	 		intermediate[4095+337:0+337] <= intermediate[4095+337:0+337] + a; end
12'd338: begin if(a[338]==1) 
	 		intermediate[4095+338:0+338] <= intermediate[4095+338:0+338] + a; end
12'd339: begin if(a[339]==1) 
	 		intermediate[4095+339:0+339] <= intermediate[4095+339:0+339] + a; end
12'd340: begin if(a[340]==1) 
	 		intermediate[4095+340:0+340] <= intermediate[4095+340:0+340] + a; end
12'd341: begin if(a[341]==1) 
	 		intermediate[4095+341:0+341] <= intermediate[4095+341:0+341] + a; end
12'd342: begin if(a[342]==1) 
	 		intermediate[4095+342:0+342] <= intermediate[4095+342:0+342] + a; end
12'd343: begin if(a[343]==1) 
	 		intermediate[4095+343:0+343] <= intermediate[4095+343:0+343] + a; end
12'd344: begin if(a[344]==1) 
	 		intermediate[4095+344:0+344] <= intermediate[4095+344:0+344] + a; end
12'd345: begin if(a[345]==1) 
	 		intermediate[4095+345:0+345] <= intermediate[4095+345:0+345] + a; end
12'd346: begin if(a[346]==1) 
	 		intermediate[4095+346:0+346] <= intermediate[4095+346:0+346] + a; end
12'd347: begin if(a[347]==1) 
	 		intermediate[4095+347:0+347] <= intermediate[4095+347:0+347] + a; end
12'd348: begin if(a[348]==1) 
	 		intermediate[4095+348:0+348] <= intermediate[4095+348:0+348] + a; end
12'd349: begin if(a[349]==1) 
	 		intermediate[4095+349:0+349] <= intermediate[4095+349:0+349] + a; end
12'd350: begin if(a[350]==1) 
	 		intermediate[4095+350:0+350] <= intermediate[4095+350:0+350] + a; end
12'd351: begin if(a[351]==1) 
	 		intermediate[4095+351:0+351] <= intermediate[4095+351:0+351] + a; end
12'd352: begin if(a[352]==1) 
	 		intermediate[4095+352:0+352] <= intermediate[4095+352:0+352] + a; end
12'd353: begin if(a[353]==1) 
	 		intermediate[4095+353:0+353] <= intermediate[4095+353:0+353] + a; end
12'd354: begin if(a[354]==1) 
	 		intermediate[4095+354:0+354] <= intermediate[4095+354:0+354] + a; end
12'd355: begin if(a[355]==1) 
	 		intermediate[4095+355:0+355] <= intermediate[4095+355:0+355] + a; end
12'd356: begin if(a[356]==1) 
	 		intermediate[4095+356:0+356] <= intermediate[4095+356:0+356] + a; end
12'd357: begin if(a[357]==1) 
	 		intermediate[4095+357:0+357] <= intermediate[4095+357:0+357] + a; end
12'd358: begin if(a[358]==1) 
	 		intermediate[4095+358:0+358] <= intermediate[4095+358:0+358] + a; end
12'd359: begin if(a[359]==1) 
	 		intermediate[4095+359:0+359] <= intermediate[4095+359:0+359] + a; end
12'd360: begin if(a[360]==1) 
	 		intermediate[4095+360:0+360] <= intermediate[4095+360:0+360] + a; end
12'd361: begin if(a[361]==1) 
	 		intermediate[4095+361:0+361] <= intermediate[4095+361:0+361] + a; end
12'd362: begin if(a[362]==1) 
	 		intermediate[4095+362:0+362] <= intermediate[4095+362:0+362] + a; end
12'd363: begin if(a[363]==1) 
	 		intermediate[4095+363:0+363] <= intermediate[4095+363:0+363] + a; end
12'd364: begin if(a[364]==1) 
	 		intermediate[4095+364:0+364] <= intermediate[4095+364:0+364] + a; end
12'd365: begin if(a[365]==1) 
	 		intermediate[4095+365:0+365] <= intermediate[4095+365:0+365] + a; end
12'd366: begin if(a[366]==1) 
	 		intermediate[4095+366:0+366] <= intermediate[4095+366:0+366] + a; end
12'd367: begin if(a[367]==1) 
	 		intermediate[4095+367:0+367] <= intermediate[4095+367:0+367] + a; end
12'd368: begin if(a[368]==1) 
	 		intermediate[4095+368:0+368] <= intermediate[4095+368:0+368] + a; end
12'd369: begin if(a[369]==1) 
	 		intermediate[4095+369:0+369] <= intermediate[4095+369:0+369] + a; end
12'd370: begin if(a[370]==1) 
	 		intermediate[4095+370:0+370] <= intermediate[4095+370:0+370] + a; end
12'd371: begin if(a[371]==1) 
	 		intermediate[4095+371:0+371] <= intermediate[4095+371:0+371] + a; end
12'd372: begin if(a[372]==1) 
	 		intermediate[4095+372:0+372] <= intermediate[4095+372:0+372] + a; end
12'd373: begin if(a[373]==1) 
	 		intermediate[4095+373:0+373] <= intermediate[4095+373:0+373] + a; end
12'd374: begin if(a[374]==1) 
	 		intermediate[4095+374:0+374] <= intermediate[4095+374:0+374] + a; end
12'd375: begin if(a[375]==1) 
	 		intermediate[4095+375:0+375] <= intermediate[4095+375:0+375] + a; end
12'd376: begin if(a[376]==1) 
	 		intermediate[4095+376:0+376] <= intermediate[4095+376:0+376] + a; end
12'd377: begin if(a[377]==1) 
	 		intermediate[4095+377:0+377] <= intermediate[4095+377:0+377] + a; end
12'd378: begin if(a[378]==1) 
	 		intermediate[4095+378:0+378] <= intermediate[4095+378:0+378] + a; end
12'd379: begin if(a[379]==1) 
	 		intermediate[4095+379:0+379] <= intermediate[4095+379:0+379] + a; end
12'd380: begin if(a[380]==1) 
	 		intermediate[4095+380:0+380] <= intermediate[4095+380:0+380] + a; end
12'd381: begin if(a[381]==1) 
	 		intermediate[4095+381:0+381] <= intermediate[4095+381:0+381] + a; end
12'd382: begin if(a[382]==1) 
	 		intermediate[4095+382:0+382] <= intermediate[4095+382:0+382] + a; end
12'd383: begin if(a[383]==1) 
	 		intermediate[4095+383:0+383] <= intermediate[4095+383:0+383] + a; end
12'd384: begin if(a[384]==1) 
	 		intermediate[4095+384:0+384] <= intermediate[4095+384:0+384] + a; end
12'd385: begin if(a[385]==1) 
	 		intermediate[4095+385:0+385] <= intermediate[4095+385:0+385] + a; end
12'd386: begin if(a[386]==1) 
	 		intermediate[4095+386:0+386] <= intermediate[4095+386:0+386] + a; end
12'd387: begin if(a[387]==1) 
	 		intermediate[4095+387:0+387] <= intermediate[4095+387:0+387] + a; end
12'd388: begin if(a[388]==1) 
	 		intermediate[4095+388:0+388] <= intermediate[4095+388:0+388] + a; end
12'd389: begin if(a[389]==1) 
	 		intermediate[4095+389:0+389] <= intermediate[4095+389:0+389] + a; end
12'd390: begin if(a[390]==1) 
	 		intermediate[4095+390:0+390] <= intermediate[4095+390:0+390] + a; end
12'd391: begin if(a[391]==1) 
	 		intermediate[4095+391:0+391] <= intermediate[4095+391:0+391] + a; end
12'd392: begin if(a[392]==1) 
	 		intermediate[4095+392:0+392] <= intermediate[4095+392:0+392] + a; end
12'd393: begin if(a[393]==1) 
	 		intermediate[4095+393:0+393] <= intermediate[4095+393:0+393] + a; end
12'd394: begin if(a[394]==1) 
	 		intermediate[4095+394:0+394] <= intermediate[4095+394:0+394] + a; end
12'd395: begin if(a[395]==1) 
	 		intermediate[4095+395:0+395] <= intermediate[4095+395:0+395] + a; end
12'd396: begin if(a[396]==1) 
	 		intermediate[4095+396:0+396] <= intermediate[4095+396:0+396] + a; end
12'd397: begin if(a[397]==1) 
	 		intermediate[4095+397:0+397] <= intermediate[4095+397:0+397] + a; end
12'd398: begin if(a[398]==1) 
	 		intermediate[4095+398:0+398] <= intermediate[4095+398:0+398] + a; end
12'd399: begin if(a[399]==1) 
	 		intermediate[4095+399:0+399] <= intermediate[4095+399:0+399] + a; end
12'd400: begin if(a[400]==1) 
	 		intermediate[4095+400:0+400] <= intermediate[4095+400:0+400] + a; end
12'd401: begin if(a[401]==1) 
	 		intermediate[4095+401:0+401] <= intermediate[4095+401:0+401] + a; end
12'd402: begin if(a[402]==1) 
	 		intermediate[4095+402:0+402] <= intermediate[4095+402:0+402] + a; end
12'd403: begin if(a[403]==1) 
	 		intermediate[4095+403:0+403] <= intermediate[4095+403:0+403] + a; end
12'd404: begin if(a[404]==1) 
	 		intermediate[4095+404:0+404] <= intermediate[4095+404:0+404] + a; end
12'd405: begin if(a[405]==1) 
	 		intermediate[4095+405:0+405] <= intermediate[4095+405:0+405] + a; end
12'd406: begin if(a[406]==1) 
	 		intermediate[4095+406:0+406] <= intermediate[4095+406:0+406] + a; end
12'd407: begin if(a[407]==1) 
	 		intermediate[4095+407:0+407] <= intermediate[4095+407:0+407] + a; end
12'd408: begin if(a[408]==1) 
	 		intermediate[4095+408:0+408] <= intermediate[4095+408:0+408] + a; end
12'd409: begin if(a[409]==1) 
	 		intermediate[4095+409:0+409] <= intermediate[4095+409:0+409] + a; end
12'd410: begin if(a[410]==1) 
	 		intermediate[4095+410:0+410] <= intermediate[4095+410:0+410] + a; end
12'd411: begin if(a[411]==1) 
	 		intermediate[4095+411:0+411] <= intermediate[4095+411:0+411] + a; end
12'd412: begin if(a[412]==1) 
	 		intermediate[4095+412:0+412] <= intermediate[4095+412:0+412] + a; end
12'd413: begin if(a[413]==1) 
	 		intermediate[4095+413:0+413] <= intermediate[4095+413:0+413] + a; end
12'd414: begin if(a[414]==1) 
	 		intermediate[4095+414:0+414] <= intermediate[4095+414:0+414] + a; end
12'd415: begin if(a[415]==1) 
	 		intermediate[4095+415:0+415] <= intermediate[4095+415:0+415] + a; end
12'd416: begin if(a[416]==1) 
	 		intermediate[4095+416:0+416] <= intermediate[4095+416:0+416] + a; end
12'd417: begin if(a[417]==1) 
	 		intermediate[4095+417:0+417] <= intermediate[4095+417:0+417] + a; end
12'd418: begin if(a[418]==1) 
	 		intermediate[4095+418:0+418] <= intermediate[4095+418:0+418] + a; end
12'd419: begin if(a[419]==1) 
	 		intermediate[4095+419:0+419] <= intermediate[4095+419:0+419] + a; end
12'd420: begin if(a[420]==1) 
	 		intermediate[4095+420:0+420] <= intermediate[4095+420:0+420] + a; end
12'd421: begin if(a[421]==1) 
	 		intermediate[4095+421:0+421] <= intermediate[4095+421:0+421] + a; end
12'd422: begin if(a[422]==1) 
	 		intermediate[4095+422:0+422] <= intermediate[4095+422:0+422] + a; end
12'd423: begin if(a[423]==1) 
	 		intermediate[4095+423:0+423] <= intermediate[4095+423:0+423] + a; end
12'd424: begin if(a[424]==1) 
	 		intermediate[4095+424:0+424] <= intermediate[4095+424:0+424] + a; end
12'd425: begin if(a[425]==1) 
	 		intermediate[4095+425:0+425] <= intermediate[4095+425:0+425] + a; end
12'd426: begin if(a[426]==1) 
	 		intermediate[4095+426:0+426] <= intermediate[4095+426:0+426] + a; end
12'd427: begin if(a[427]==1) 
	 		intermediate[4095+427:0+427] <= intermediate[4095+427:0+427] + a; end
12'd428: begin if(a[428]==1) 
	 		intermediate[4095+428:0+428] <= intermediate[4095+428:0+428] + a; end
12'd429: begin if(a[429]==1) 
	 		intermediate[4095+429:0+429] <= intermediate[4095+429:0+429] + a; end
12'd430: begin if(a[430]==1) 
	 		intermediate[4095+430:0+430] <= intermediate[4095+430:0+430] + a; end
12'd431: begin if(a[431]==1) 
	 		intermediate[4095+431:0+431] <= intermediate[4095+431:0+431] + a; end
12'd432: begin if(a[432]==1) 
	 		intermediate[4095+432:0+432] <= intermediate[4095+432:0+432] + a; end
12'd433: begin if(a[433]==1) 
	 		intermediate[4095+433:0+433] <= intermediate[4095+433:0+433] + a; end
12'd434: begin if(a[434]==1) 
	 		intermediate[4095+434:0+434] <= intermediate[4095+434:0+434] + a; end
12'd435: begin if(a[435]==1) 
	 		intermediate[4095+435:0+435] <= intermediate[4095+435:0+435] + a; end
12'd436: begin if(a[436]==1) 
	 		intermediate[4095+436:0+436] <= intermediate[4095+436:0+436] + a; end
12'd437: begin if(a[437]==1) 
	 		intermediate[4095+437:0+437] <= intermediate[4095+437:0+437] + a; end
12'd438: begin if(a[438]==1) 
	 		intermediate[4095+438:0+438] <= intermediate[4095+438:0+438] + a; end
12'd439: begin if(a[439]==1) 
	 		intermediate[4095+439:0+439] <= intermediate[4095+439:0+439] + a; end
12'd440: begin if(a[440]==1) 
	 		intermediate[4095+440:0+440] <= intermediate[4095+440:0+440] + a; end
12'd441: begin if(a[441]==1) 
	 		intermediate[4095+441:0+441] <= intermediate[4095+441:0+441] + a; end
12'd442: begin if(a[442]==1) 
	 		intermediate[4095+442:0+442] <= intermediate[4095+442:0+442] + a; end
12'd443: begin if(a[443]==1) 
	 		intermediate[4095+443:0+443] <= intermediate[4095+443:0+443] + a; end
12'd444: begin if(a[444]==1) 
	 		intermediate[4095+444:0+444] <= intermediate[4095+444:0+444] + a; end
12'd445: begin if(a[445]==1) 
	 		intermediate[4095+445:0+445] <= intermediate[4095+445:0+445] + a; end
12'd446: begin if(a[446]==1) 
	 		intermediate[4095+446:0+446] <= intermediate[4095+446:0+446] + a; end
12'd447: begin if(a[447]==1) 
	 		intermediate[4095+447:0+447] <= intermediate[4095+447:0+447] + a; end
12'd448: begin if(a[448]==1) 
	 		intermediate[4095+448:0+448] <= intermediate[4095+448:0+448] + a; end
12'd449: begin if(a[449]==1) 
	 		intermediate[4095+449:0+449] <= intermediate[4095+449:0+449] + a; end
12'd450: begin if(a[450]==1) 
	 		intermediate[4095+450:0+450] <= intermediate[4095+450:0+450] + a; end
12'd451: begin if(a[451]==1) 
	 		intermediate[4095+451:0+451] <= intermediate[4095+451:0+451] + a; end
12'd452: begin if(a[452]==1) 
	 		intermediate[4095+452:0+452] <= intermediate[4095+452:0+452] + a; end
12'd453: begin if(a[453]==1) 
	 		intermediate[4095+453:0+453] <= intermediate[4095+453:0+453] + a; end
12'd454: begin if(a[454]==1) 
	 		intermediate[4095+454:0+454] <= intermediate[4095+454:0+454] + a; end
12'd455: begin if(a[455]==1) 
	 		intermediate[4095+455:0+455] <= intermediate[4095+455:0+455] + a; end
12'd456: begin if(a[456]==1) 
	 		intermediate[4095+456:0+456] <= intermediate[4095+456:0+456] + a; end
12'd457: begin if(a[457]==1) 
	 		intermediate[4095+457:0+457] <= intermediate[4095+457:0+457] + a; end
12'd458: begin if(a[458]==1) 
	 		intermediate[4095+458:0+458] <= intermediate[4095+458:0+458] + a; end
12'd459: begin if(a[459]==1) 
	 		intermediate[4095+459:0+459] <= intermediate[4095+459:0+459] + a; end
12'd460: begin if(a[460]==1) 
	 		intermediate[4095+460:0+460] <= intermediate[4095+460:0+460] + a; end
12'd461: begin if(a[461]==1) 
	 		intermediate[4095+461:0+461] <= intermediate[4095+461:0+461] + a; end
12'd462: begin if(a[462]==1) 
	 		intermediate[4095+462:0+462] <= intermediate[4095+462:0+462] + a; end
12'd463: begin if(a[463]==1) 
	 		intermediate[4095+463:0+463] <= intermediate[4095+463:0+463] + a; end
12'd464: begin if(a[464]==1) 
	 		intermediate[4095+464:0+464] <= intermediate[4095+464:0+464] + a; end
12'd465: begin if(a[465]==1) 
	 		intermediate[4095+465:0+465] <= intermediate[4095+465:0+465] + a; end
12'd466: begin if(a[466]==1) 
	 		intermediate[4095+466:0+466] <= intermediate[4095+466:0+466] + a; end
12'd467: begin if(a[467]==1) 
	 		intermediate[4095+467:0+467] <= intermediate[4095+467:0+467] + a; end
12'd468: begin if(a[468]==1) 
	 		intermediate[4095+468:0+468] <= intermediate[4095+468:0+468] + a; end
12'd469: begin if(a[469]==1) 
	 		intermediate[4095+469:0+469] <= intermediate[4095+469:0+469] + a; end
12'd470: begin if(a[470]==1) 
	 		intermediate[4095+470:0+470] <= intermediate[4095+470:0+470] + a; end
12'd471: begin if(a[471]==1) 
	 		intermediate[4095+471:0+471] <= intermediate[4095+471:0+471] + a; end
12'd472: begin if(a[472]==1) 
	 		intermediate[4095+472:0+472] <= intermediate[4095+472:0+472] + a; end
12'd473: begin if(a[473]==1) 
	 		intermediate[4095+473:0+473] <= intermediate[4095+473:0+473] + a; end
12'd474: begin if(a[474]==1) 
	 		intermediate[4095+474:0+474] <= intermediate[4095+474:0+474] + a; end
12'd475: begin if(a[475]==1) 
	 		intermediate[4095+475:0+475] <= intermediate[4095+475:0+475] + a; end
12'd476: begin if(a[476]==1) 
	 		intermediate[4095+476:0+476] <= intermediate[4095+476:0+476] + a; end
12'd477: begin if(a[477]==1) 
	 		intermediate[4095+477:0+477] <= intermediate[4095+477:0+477] + a; end
12'd478: begin if(a[478]==1) 
	 		intermediate[4095+478:0+478] <= intermediate[4095+478:0+478] + a; end
12'd479: begin if(a[479]==1) 
	 		intermediate[4095+479:0+479] <= intermediate[4095+479:0+479] + a; end
12'd480: begin if(a[480]==1) 
	 		intermediate[4095+480:0+480] <= intermediate[4095+480:0+480] + a; end
12'd481: begin if(a[481]==1) 
	 		intermediate[4095+481:0+481] <= intermediate[4095+481:0+481] + a; end
12'd482: begin if(a[482]==1) 
	 		intermediate[4095+482:0+482] <= intermediate[4095+482:0+482] + a; end
12'd483: begin if(a[483]==1) 
	 		intermediate[4095+483:0+483] <= intermediate[4095+483:0+483] + a; end
12'd484: begin if(a[484]==1) 
	 		intermediate[4095+484:0+484] <= intermediate[4095+484:0+484] + a; end
12'd485: begin if(a[485]==1) 
	 		intermediate[4095+485:0+485] <= intermediate[4095+485:0+485] + a; end
12'd486: begin if(a[486]==1) 
	 		intermediate[4095+486:0+486] <= intermediate[4095+486:0+486] + a; end
12'd487: begin if(a[487]==1) 
	 		intermediate[4095+487:0+487] <= intermediate[4095+487:0+487] + a; end
12'd488: begin if(a[488]==1) 
	 		intermediate[4095+488:0+488] <= intermediate[4095+488:0+488] + a; end
12'd489: begin if(a[489]==1) 
	 		intermediate[4095+489:0+489] <= intermediate[4095+489:0+489] + a; end
12'd490: begin if(a[490]==1) 
	 		intermediate[4095+490:0+490] <= intermediate[4095+490:0+490] + a; end
12'd491: begin if(a[491]==1) 
	 		intermediate[4095+491:0+491] <= intermediate[4095+491:0+491] + a; end
12'd492: begin if(a[492]==1) 
	 		intermediate[4095+492:0+492] <= intermediate[4095+492:0+492] + a; end
12'd493: begin if(a[493]==1) 
	 		intermediate[4095+493:0+493] <= intermediate[4095+493:0+493] + a; end
12'd494: begin if(a[494]==1) 
	 		intermediate[4095+494:0+494] <= intermediate[4095+494:0+494] + a; end
12'd495: begin if(a[495]==1) 
	 		intermediate[4095+495:0+495] <= intermediate[4095+495:0+495] + a; end
12'd496: begin if(a[496]==1) 
	 		intermediate[4095+496:0+496] <= intermediate[4095+496:0+496] + a; end
12'd497: begin if(a[497]==1) 
	 		intermediate[4095+497:0+497] <= intermediate[4095+497:0+497] + a; end
12'd498: begin if(a[498]==1) 
	 		intermediate[4095+498:0+498] <= intermediate[4095+498:0+498] + a; end
12'd499: begin if(a[499]==1) 
	 		intermediate[4095+499:0+499] <= intermediate[4095+499:0+499] + a; end
12'd500: begin if(a[500]==1) 
	 		intermediate[4095+500:0+500] <= intermediate[4095+500:0+500] + a; end
12'd501: begin if(a[501]==1) 
	 		intermediate[4095+501:0+501] <= intermediate[4095+501:0+501] + a; end
12'd502: begin if(a[502]==1) 
	 		intermediate[4095+502:0+502] <= intermediate[4095+502:0+502] + a; end
12'd503: begin if(a[503]==1) 
	 		intermediate[4095+503:0+503] <= intermediate[4095+503:0+503] + a; end
12'd504: begin if(a[504]==1) 
	 		intermediate[4095+504:0+504] <= intermediate[4095+504:0+504] + a; end
12'd505: begin if(a[505]==1) 
	 		intermediate[4095+505:0+505] <= intermediate[4095+505:0+505] + a; end
12'd506: begin if(a[506]==1) 
	 		intermediate[4095+506:0+506] <= intermediate[4095+506:0+506] + a; end
12'd507: begin if(a[507]==1) 
	 		intermediate[4095+507:0+507] <= intermediate[4095+507:0+507] + a; end
12'd508: begin if(a[508]==1) 
	 		intermediate[4095+508:0+508] <= intermediate[4095+508:0+508] + a; end
12'd509: begin if(a[509]==1) 
	 		intermediate[4095+509:0+509] <= intermediate[4095+509:0+509] + a; end
12'd510: begin if(a[510]==1) 
	 		intermediate[4095+510:0+510] <= intermediate[4095+510:0+510] + a; end
12'd511: begin if(a[511]==1) 
	 		intermediate[4095+511:0+511] <= intermediate[4095+511:0+511] + a; end
12'd512: begin if(a[512]==1) 
	 		intermediate[4095+512:0+512] <= intermediate[4095+512:0+512] + a; end
12'd513: begin if(a[513]==1) 
	 		intermediate[4095+513:0+513] <= intermediate[4095+513:0+513] + a; end
12'd514: begin if(a[514]==1) 
	 		intermediate[4095+514:0+514] <= intermediate[4095+514:0+514] + a; end
12'd515: begin if(a[515]==1) 
	 		intermediate[4095+515:0+515] <= intermediate[4095+515:0+515] + a; end
12'd516: begin if(a[516]==1) 
	 		intermediate[4095+516:0+516] <= intermediate[4095+516:0+516] + a; end
12'd517: begin if(a[517]==1) 
	 		intermediate[4095+517:0+517] <= intermediate[4095+517:0+517] + a; end
12'd518: begin if(a[518]==1) 
	 		intermediate[4095+518:0+518] <= intermediate[4095+518:0+518] + a; end
12'd519: begin if(a[519]==1) 
	 		intermediate[4095+519:0+519] <= intermediate[4095+519:0+519] + a; end
12'd520: begin if(a[520]==1) 
	 		intermediate[4095+520:0+520] <= intermediate[4095+520:0+520] + a; end
12'd521: begin if(a[521]==1) 
	 		intermediate[4095+521:0+521] <= intermediate[4095+521:0+521] + a; end
12'd522: begin if(a[522]==1) 
	 		intermediate[4095+522:0+522] <= intermediate[4095+522:0+522] + a; end
12'd523: begin if(a[523]==1) 
	 		intermediate[4095+523:0+523] <= intermediate[4095+523:0+523] + a; end
12'd524: begin if(a[524]==1) 
	 		intermediate[4095+524:0+524] <= intermediate[4095+524:0+524] + a; end
12'd525: begin if(a[525]==1) 
	 		intermediate[4095+525:0+525] <= intermediate[4095+525:0+525] + a; end
12'd526: begin if(a[526]==1) 
	 		intermediate[4095+526:0+526] <= intermediate[4095+526:0+526] + a; end
12'd527: begin if(a[527]==1) 
	 		intermediate[4095+527:0+527] <= intermediate[4095+527:0+527] + a; end
12'd528: begin if(a[528]==1) 
	 		intermediate[4095+528:0+528] <= intermediate[4095+528:0+528] + a; end
12'd529: begin if(a[529]==1) 
	 		intermediate[4095+529:0+529] <= intermediate[4095+529:0+529] + a; end
12'd530: begin if(a[530]==1) 
	 		intermediate[4095+530:0+530] <= intermediate[4095+530:0+530] + a; end
12'd531: begin if(a[531]==1) 
	 		intermediate[4095+531:0+531] <= intermediate[4095+531:0+531] + a; end
12'd532: begin if(a[532]==1) 
	 		intermediate[4095+532:0+532] <= intermediate[4095+532:0+532] + a; end
12'd533: begin if(a[533]==1) 
	 		intermediate[4095+533:0+533] <= intermediate[4095+533:0+533] + a; end
12'd534: begin if(a[534]==1) 
	 		intermediate[4095+534:0+534] <= intermediate[4095+534:0+534] + a; end
12'd535: begin if(a[535]==1) 
	 		intermediate[4095+535:0+535] <= intermediate[4095+535:0+535] + a; end
12'd536: begin if(a[536]==1) 
	 		intermediate[4095+536:0+536] <= intermediate[4095+536:0+536] + a; end
12'd537: begin if(a[537]==1) 
	 		intermediate[4095+537:0+537] <= intermediate[4095+537:0+537] + a; end
12'd538: begin if(a[538]==1) 
	 		intermediate[4095+538:0+538] <= intermediate[4095+538:0+538] + a; end
12'd539: begin if(a[539]==1) 
	 		intermediate[4095+539:0+539] <= intermediate[4095+539:0+539] + a; end
12'd540: begin if(a[540]==1) 
	 		intermediate[4095+540:0+540] <= intermediate[4095+540:0+540] + a; end
12'd541: begin if(a[541]==1) 
	 		intermediate[4095+541:0+541] <= intermediate[4095+541:0+541] + a; end
12'd542: begin if(a[542]==1) 
	 		intermediate[4095+542:0+542] <= intermediate[4095+542:0+542] + a; end
12'd543: begin if(a[543]==1) 
	 		intermediate[4095+543:0+543] <= intermediate[4095+543:0+543] + a; end
12'd544: begin if(a[544]==1) 
	 		intermediate[4095+544:0+544] <= intermediate[4095+544:0+544] + a; end
12'd545: begin if(a[545]==1) 
	 		intermediate[4095+545:0+545] <= intermediate[4095+545:0+545] + a; end
12'd546: begin if(a[546]==1) 
	 		intermediate[4095+546:0+546] <= intermediate[4095+546:0+546] + a; end
12'd547: begin if(a[547]==1) 
	 		intermediate[4095+547:0+547] <= intermediate[4095+547:0+547] + a; end
12'd548: begin if(a[548]==1) 
	 		intermediate[4095+548:0+548] <= intermediate[4095+548:0+548] + a; end
12'd549: begin if(a[549]==1) 
	 		intermediate[4095+549:0+549] <= intermediate[4095+549:0+549] + a; end
12'd550: begin if(a[550]==1) 
	 		intermediate[4095+550:0+550] <= intermediate[4095+550:0+550] + a; end
12'd551: begin if(a[551]==1) 
	 		intermediate[4095+551:0+551] <= intermediate[4095+551:0+551] + a; end
12'd552: begin if(a[552]==1) 
	 		intermediate[4095+552:0+552] <= intermediate[4095+552:0+552] + a; end
12'd553: begin if(a[553]==1) 
	 		intermediate[4095+553:0+553] <= intermediate[4095+553:0+553] + a; end
12'd554: begin if(a[554]==1) 
	 		intermediate[4095+554:0+554] <= intermediate[4095+554:0+554] + a; end
12'd555: begin if(a[555]==1) 
	 		intermediate[4095+555:0+555] <= intermediate[4095+555:0+555] + a; end
12'd556: begin if(a[556]==1) 
	 		intermediate[4095+556:0+556] <= intermediate[4095+556:0+556] + a; end
12'd557: begin if(a[557]==1) 
	 		intermediate[4095+557:0+557] <= intermediate[4095+557:0+557] + a; end
12'd558: begin if(a[558]==1) 
	 		intermediate[4095+558:0+558] <= intermediate[4095+558:0+558] + a; end
12'd559: begin if(a[559]==1) 
	 		intermediate[4095+559:0+559] <= intermediate[4095+559:0+559] + a; end
12'd560: begin if(a[560]==1) 
	 		intermediate[4095+560:0+560] <= intermediate[4095+560:0+560] + a; end
12'd561: begin if(a[561]==1) 
	 		intermediate[4095+561:0+561] <= intermediate[4095+561:0+561] + a; end
12'd562: begin if(a[562]==1) 
	 		intermediate[4095+562:0+562] <= intermediate[4095+562:0+562] + a; end
12'd563: begin if(a[563]==1) 
	 		intermediate[4095+563:0+563] <= intermediate[4095+563:0+563] + a; end
12'd564: begin if(a[564]==1) 
	 		intermediate[4095+564:0+564] <= intermediate[4095+564:0+564] + a; end
12'd565: begin if(a[565]==1) 
	 		intermediate[4095+565:0+565] <= intermediate[4095+565:0+565] + a; end
12'd566: begin if(a[566]==1) 
	 		intermediate[4095+566:0+566] <= intermediate[4095+566:0+566] + a; end
12'd567: begin if(a[567]==1) 
	 		intermediate[4095+567:0+567] <= intermediate[4095+567:0+567] + a; end
12'd568: begin if(a[568]==1) 
	 		intermediate[4095+568:0+568] <= intermediate[4095+568:0+568] + a; end
12'd569: begin if(a[569]==1) 
	 		intermediate[4095+569:0+569] <= intermediate[4095+569:0+569] + a; end
12'd570: begin if(a[570]==1) 
	 		intermediate[4095+570:0+570] <= intermediate[4095+570:0+570] + a; end
12'd571: begin if(a[571]==1) 
	 		intermediate[4095+571:0+571] <= intermediate[4095+571:0+571] + a; end
12'd572: begin if(a[572]==1) 
	 		intermediate[4095+572:0+572] <= intermediate[4095+572:0+572] + a; end
12'd573: begin if(a[573]==1) 
	 		intermediate[4095+573:0+573] <= intermediate[4095+573:0+573] + a; end
12'd574: begin if(a[574]==1) 
	 		intermediate[4095+574:0+574] <= intermediate[4095+574:0+574] + a; end
12'd575: begin if(a[575]==1) 
	 		intermediate[4095+575:0+575] <= intermediate[4095+575:0+575] + a; end
12'd576: begin if(a[576]==1) 
	 		intermediate[4095+576:0+576] <= intermediate[4095+576:0+576] + a; end
12'd577: begin if(a[577]==1) 
	 		intermediate[4095+577:0+577] <= intermediate[4095+577:0+577] + a; end
12'd578: begin if(a[578]==1) 
	 		intermediate[4095+578:0+578] <= intermediate[4095+578:0+578] + a; end
12'd579: begin if(a[579]==1) 
	 		intermediate[4095+579:0+579] <= intermediate[4095+579:0+579] + a; end
12'd580: begin if(a[580]==1) 
	 		intermediate[4095+580:0+580] <= intermediate[4095+580:0+580] + a; end
12'd581: begin if(a[581]==1) 
	 		intermediate[4095+581:0+581] <= intermediate[4095+581:0+581] + a; end
12'd582: begin if(a[582]==1) 
	 		intermediate[4095+582:0+582] <= intermediate[4095+582:0+582] + a; end
12'd583: begin if(a[583]==1) 
	 		intermediate[4095+583:0+583] <= intermediate[4095+583:0+583] + a; end
12'd584: begin if(a[584]==1) 
	 		intermediate[4095+584:0+584] <= intermediate[4095+584:0+584] + a; end
12'd585: begin if(a[585]==1) 
	 		intermediate[4095+585:0+585] <= intermediate[4095+585:0+585] + a; end
12'd586: begin if(a[586]==1) 
	 		intermediate[4095+586:0+586] <= intermediate[4095+586:0+586] + a; end
12'd587: begin if(a[587]==1) 
	 		intermediate[4095+587:0+587] <= intermediate[4095+587:0+587] + a; end
12'd588: begin if(a[588]==1) 
	 		intermediate[4095+588:0+588] <= intermediate[4095+588:0+588] + a; end
12'd589: begin if(a[589]==1) 
	 		intermediate[4095+589:0+589] <= intermediate[4095+589:0+589] + a; end
12'd590: begin if(a[590]==1) 
	 		intermediate[4095+590:0+590] <= intermediate[4095+590:0+590] + a; end
12'd591: begin if(a[591]==1) 
	 		intermediate[4095+591:0+591] <= intermediate[4095+591:0+591] + a; end
12'd592: begin if(a[592]==1) 
	 		intermediate[4095+592:0+592] <= intermediate[4095+592:0+592] + a; end
12'd593: begin if(a[593]==1) 
	 		intermediate[4095+593:0+593] <= intermediate[4095+593:0+593] + a; end
12'd594: begin if(a[594]==1) 
	 		intermediate[4095+594:0+594] <= intermediate[4095+594:0+594] + a; end
12'd595: begin if(a[595]==1) 
	 		intermediate[4095+595:0+595] <= intermediate[4095+595:0+595] + a; end
12'd596: begin if(a[596]==1) 
	 		intermediate[4095+596:0+596] <= intermediate[4095+596:0+596] + a; end
12'd597: begin if(a[597]==1) 
	 		intermediate[4095+597:0+597] <= intermediate[4095+597:0+597] + a; end
12'd598: begin if(a[598]==1) 
	 		intermediate[4095+598:0+598] <= intermediate[4095+598:0+598] + a; end
12'd599: begin if(a[599]==1) 
	 		intermediate[4095+599:0+599] <= intermediate[4095+599:0+599] + a; end
12'd600: begin if(a[600]==1) 
	 		intermediate[4095+600:0+600] <= intermediate[4095+600:0+600] + a; end
12'd601: begin if(a[601]==1) 
	 		intermediate[4095+601:0+601] <= intermediate[4095+601:0+601] + a; end
12'd602: begin if(a[602]==1) 
	 		intermediate[4095+602:0+602] <= intermediate[4095+602:0+602] + a; end
12'd603: begin if(a[603]==1) 
	 		intermediate[4095+603:0+603] <= intermediate[4095+603:0+603] + a; end
12'd604: begin if(a[604]==1) 
	 		intermediate[4095+604:0+604] <= intermediate[4095+604:0+604] + a; end
12'd605: begin if(a[605]==1) 
	 		intermediate[4095+605:0+605] <= intermediate[4095+605:0+605] + a; end
12'd606: begin if(a[606]==1) 
	 		intermediate[4095+606:0+606] <= intermediate[4095+606:0+606] + a; end
12'd607: begin if(a[607]==1) 
	 		intermediate[4095+607:0+607] <= intermediate[4095+607:0+607] + a; end
12'd608: begin if(a[608]==1) 
	 		intermediate[4095+608:0+608] <= intermediate[4095+608:0+608] + a; end
12'd609: begin if(a[609]==1) 
	 		intermediate[4095+609:0+609] <= intermediate[4095+609:0+609] + a; end
12'd610: begin if(a[610]==1) 
	 		intermediate[4095+610:0+610] <= intermediate[4095+610:0+610] + a; end
12'd611: begin if(a[611]==1) 
	 		intermediate[4095+611:0+611] <= intermediate[4095+611:0+611] + a; end
12'd612: begin if(a[612]==1) 
	 		intermediate[4095+612:0+612] <= intermediate[4095+612:0+612] + a; end
12'd613: begin if(a[613]==1) 
	 		intermediate[4095+613:0+613] <= intermediate[4095+613:0+613] + a; end
12'd614: begin if(a[614]==1) 
	 		intermediate[4095+614:0+614] <= intermediate[4095+614:0+614] + a; end
12'd615: begin if(a[615]==1) 
	 		intermediate[4095+615:0+615] <= intermediate[4095+615:0+615] + a; end
12'd616: begin if(a[616]==1) 
	 		intermediate[4095+616:0+616] <= intermediate[4095+616:0+616] + a; end
12'd617: begin if(a[617]==1) 
	 		intermediate[4095+617:0+617] <= intermediate[4095+617:0+617] + a; end
12'd618: begin if(a[618]==1) 
	 		intermediate[4095+618:0+618] <= intermediate[4095+618:0+618] + a; end
12'd619: begin if(a[619]==1) 
	 		intermediate[4095+619:0+619] <= intermediate[4095+619:0+619] + a; end
12'd620: begin if(a[620]==1) 
	 		intermediate[4095+620:0+620] <= intermediate[4095+620:0+620] + a; end
12'd621: begin if(a[621]==1) 
	 		intermediate[4095+621:0+621] <= intermediate[4095+621:0+621] + a; end
12'd622: begin if(a[622]==1) 
	 		intermediate[4095+622:0+622] <= intermediate[4095+622:0+622] + a; end
12'd623: begin if(a[623]==1) 
	 		intermediate[4095+623:0+623] <= intermediate[4095+623:0+623] + a; end
12'd624: begin if(a[624]==1) 
	 		intermediate[4095+624:0+624] <= intermediate[4095+624:0+624] + a; end
12'd625: begin if(a[625]==1) 
	 		intermediate[4095+625:0+625] <= intermediate[4095+625:0+625] + a; end
12'd626: begin if(a[626]==1) 
	 		intermediate[4095+626:0+626] <= intermediate[4095+626:0+626] + a; end
12'd627: begin if(a[627]==1) 
	 		intermediate[4095+627:0+627] <= intermediate[4095+627:0+627] + a; end
12'd628: begin if(a[628]==1) 
	 		intermediate[4095+628:0+628] <= intermediate[4095+628:0+628] + a; end
12'd629: begin if(a[629]==1) 
	 		intermediate[4095+629:0+629] <= intermediate[4095+629:0+629] + a; end
12'd630: begin if(a[630]==1) 
	 		intermediate[4095+630:0+630] <= intermediate[4095+630:0+630] + a; end
12'd631: begin if(a[631]==1) 
	 		intermediate[4095+631:0+631] <= intermediate[4095+631:0+631] + a; end
12'd632: begin if(a[632]==1) 
	 		intermediate[4095+632:0+632] <= intermediate[4095+632:0+632] + a; end
12'd633: begin if(a[633]==1) 
	 		intermediate[4095+633:0+633] <= intermediate[4095+633:0+633] + a; end
12'd634: begin if(a[634]==1) 
	 		intermediate[4095+634:0+634] <= intermediate[4095+634:0+634] + a; end
12'd635: begin if(a[635]==1) 
	 		intermediate[4095+635:0+635] <= intermediate[4095+635:0+635] + a; end
12'd636: begin if(a[636]==1) 
	 		intermediate[4095+636:0+636] <= intermediate[4095+636:0+636] + a; end
12'd637: begin if(a[637]==1) 
	 		intermediate[4095+637:0+637] <= intermediate[4095+637:0+637] + a; end
12'd638: begin if(a[638]==1) 
	 		intermediate[4095+638:0+638] <= intermediate[4095+638:0+638] + a; end
12'd639: begin if(a[639]==1) 
	 		intermediate[4095+639:0+639] <= intermediate[4095+639:0+639] + a; end
12'd640: begin if(a[640]==1) 
	 		intermediate[4095+640:0+640] <= intermediate[4095+640:0+640] + a; end
12'd641: begin if(a[641]==1) 
	 		intermediate[4095+641:0+641] <= intermediate[4095+641:0+641] + a; end
12'd642: begin if(a[642]==1) 
	 		intermediate[4095+642:0+642] <= intermediate[4095+642:0+642] + a; end
12'd643: begin if(a[643]==1) 
	 		intermediate[4095+643:0+643] <= intermediate[4095+643:0+643] + a; end
12'd644: begin if(a[644]==1) 
	 		intermediate[4095+644:0+644] <= intermediate[4095+644:0+644] + a; end
12'd645: begin if(a[645]==1) 
	 		intermediate[4095+645:0+645] <= intermediate[4095+645:0+645] + a; end
12'd646: begin if(a[646]==1) 
	 		intermediate[4095+646:0+646] <= intermediate[4095+646:0+646] + a; end
12'd647: begin if(a[647]==1) 
	 		intermediate[4095+647:0+647] <= intermediate[4095+647:0+647] + a; end
12'd648: begin if(a[648]==1) 
	 		intermediate[4095+648:0+648] <= intermediate[4095+648:0+648] + a; end
12'd649: begin if(a[649]==1) 
	 		intermediate[4095+649:0+649] <= intermediate[4095+649:0+649] + a; end
12'd650: begin if(a[650]==1) 
	 		intermediate[4095+650:0+650] <= intermediate[4095+650:0+650] + a; end
12'd651: begin if(a[651]==1) 
	 		intermediate[4095+651:0+651] <= intermediate[4095+651:0+651] + a; end
12'd652: begin if(a[652]==1) 
	 		intermediate[4095+652:0+652] <= intermediate[4095+652:0+652] + a; end
12'd653: begin if(a[653]==1) 
	 		intermediate[4095+653:0+653] <= intermediate[4095+653:0+653] + a; end
12'd654: begin if(a[654]==1) 
	 		intermediate[4095+654:0+654] <= intermediate[4095+654:0+654] + a; end
12'd655: begin if(a[655]==1) 
	 		intermediate[4095+655:0+655] <= intermediate[4095+655:0+655] + a; end
12'd656: begin if(a[656]==1) 
	 		intermediate[4095+656:0+656] <= intermediate[4095+656:0+656] + a; end
12'd657: begin if(a[657]==1) 
	 		intermediate[4095+657:0+657] <= intermediate[4095+657:0+657] + a; end
12'd658: begin if(a[658]==1) 
	 		intermediate[4095+658:0+658] <= intermediate[4095+658:0+658] + a; end
12'd659: begin if(a[659]==1) 
	 		intermediate[4095+659:0+659] <= intermediate[4095+659:0+659] + a; end
12'd660: begin if(a[660]==1) 
	 		intermediate[4095+660:0+660] <= intermediate[4095+660:0+660] + a; end
12'd661: begin if(a[661]==1) 
	 		intermediate[4095+661:0+661] <= intermediate[4095+661:0+661] + a; end
12'd662: begin if(a[662]==1) 
	 		intermediate[4095+662:0+662] <= intermediate[4095+662:0+662] + a; end
12'd663: begin if(a[663]==1) 
	 		intermediate[4095+663:0+663] <= intermediate[4095+663:0+663] + a; end
12'd664: begin if(a[664]==1) 
	 		intermediate[4095+664:0+664] <= intermediate[4095+664:0+664] + a; end
12'd665: begin if(a[665]==1) 
	 		intermediate[4095+665:0+665] <= intermediate[4095+665:0+665] + a; end
12'd666: begin if(a[666]==1) 
	 		intermediate[4095+666:0+666] <= intermediate[4095+666:0+666] + a; end
12'd667: begin if(a[667]==1) 
	 		intermediate[4095+667:0+667] <= intermediate[4095+667:0+667] + a; end
12'd668: begin if(a[668]==1) 
	 		intermediate[4095+668:0+668] <= intermediate[4095+668:0+668] + a; end
12'd669: begin if(a[669]==1) 
	 		intermediate[4095+669:0+669] <= intermediate[4095+669:0+669] + a; end
12'd670: begin if(a[670]==1) 
	 		intermediate[4095+670:0+670] <= intermediate[4095+670:0+670] + a; end
12'd671: begin if(a[671]==1) 
	 		intermediate[4095+671:0+671] <= intermediate[4095+671:0+671] + a; end
12'd672: begin if(a[672]==1) 
	 		intermediate[4095+672:0+672] <= intermediate[4095+672:0+672] + a; end
12'd673: begin if(a[673]==1) 
	 		intermediate[4095+673:0+673] <= intermediate[4095+673:0+673] + a; end
12'd674: begin if(a[674]==1) 
	 		intermediate[4095+674:0+674] <= intermediate[4095+674:0+674] + a; end
12'd675: begin if(a[675]==1) 
	 		intermediate[4095+675:0+675] <= intermediate[4095+675:0+675] + a; end
12'd676: begin if(a[676]==1) 
	 		intermediate[4095+676:0+676] <= intermediate[4095+676:0+676] + a; end
12'd677: begin if(a[677]==1) 
	 		intermediate[4095+677:0+677] <= intermediate[4095+677:0+677] + a; end
12'd678: begin if(a[678]==1) 
	 		intermediate[4095+678:0+678] <= intermediate[4095+678:0+678] + a; end
12'd679: begin if(a[679]==1) 
	 		intermediate[4095+679:0+679] <= intermediate[4095+679:0+679] + a; end
12'd680: begin if(a[680]==1) 
	 		intermediate[4095+680:0+680] <= intermediate[4095+680:0+680] + a; end
12'd681: begin if(a[681]==1) 
	 		intermediate[4095+681:0+681] <= intermediate[4095+681:0+681] + a; end
12'd682: begin if(a[682]==1) 
	 		intermediate[4095+682:0+682] <= intermediate[4095+682:0+682] + a; end
12'd683: begin if(a[683]==1) 
	 		intermediate[4095+683:0+683] <= intermediate[4095+683:0+683] + a; end
12'd684: begin if(a[684]==1) 
	 		intermediate[4095+684:0+684] <= intermediate[4095+684:0+684] + a; end
12'd685: begin if(a[685]==1) 
	 		intermediate[4095+685:0+685] <= intermediate[4095+685:0+685] + a; end
12'd686: begin if(a[686]==1) 
	 		intermediate[4095+686:0+686] <= intermediate[4095+686:0+686] + a; end
12'd687: begin if(a[687]==1) 
	 		intermediate[4095+687:0+687] <= intermediate[4095+687:0+687] + a; end
12'd688: begin if(a[688]==1) 
	 		intermediate[4095+688:0+688] <= intermediate[4095+688:0+688] + a; end
12'd689: begin if(a[689]==1) 
	 		intermediate[4095+689:0+689] <= intermediate[4095+689:0+689] + a; end
12'd690: begin if(a[690]==1) 
	 		intermediate[4095+690:0+690] <= intermediate[4095+690:0+690] + a; end
12'd691: begin if(a[691]==1) 
	 		intermediate[4095+691:0+691] <= intermediate[4095+691:0+691] + a; end
12'd692: begin if(a[692]==1) 
	 		intermediate[4095+692:0+692] <= intermediate[4095+692:0+692] + a; end
12'd693: begin if(a[693]==1) 
	 		intermediate[4095+693:0+693] <= intermediate[4095+693:0+693] + a; end
12'd694: begin if(a[694]==1) 
	 		intermediate[4095+694:0+694] <= intermediate[4095+694:0+694] + a; end
12'd695: begin if(a[695]==1) 
	 		intermediate[4095+695:0+695] <= intermediate[4095+695:0+695] + a; end
12'd696: begin if(a[696]==1) 
	 		intermediate[4095+696:0+696] <= intermediate[4095+696:0+696] + a; end
12'd697: begin if(a[697]==1) 
	 		intermediate[4095+697:0+697] <= intermediate[4095+697:0+697] + a; end
12'd698: begin if(a[698]==1) 
	 		intermediate[4095+698:0+698] <= intermediate[4095+698:0+698] + a; end
12'd699: begin if(a[699]==1) 
	 		intermediate[4095+699:0+699] <= intermediate[4095+699:0+699] + a; end
12'd700: begin if(a[700]==1) 
	 		intermediate[4095+700:0+700] <= intermediate[4095+700:0+700] + a; end
12'd701: begin if(a[701]==1) 
	 		intermediate[4095+701:0+701] <= intermediate[4095+701:0+701] + a; end
12'd702: begin if(a[702]==1) 
	 		intermediate[4095+702:0+702] <= intermediate[4095+702:0+702] + a; end
12'd703: begin if(a[703]==1) 
	 		intermediate[4095+703:0+703] <= intermediate[4095+703:0+703] + a; end
12'd704: begin if(a[704]==1) 
	 		intermediate[4095+704:0+704] <= intermediate[4095+704:0+704] + a; end
12'd705: begin if(a[705]==1) 
	 		intermediate[4095+705:0+705] <= intermediate[4095+705:0+705] + a; end
12'd706: begin if(a[706]==1) 
	 		intermediate[4095+706:0+706] <= intermediate[4095+706:0+706] + a; end
12'd707: begin if(a[707]==1) 
	 		intermediate[4095+707:0+707] <= intermediate[4095+707:0+707] + a; end
12'd708: begin if(a[708]==1) 
	 		intermediate[4095+708:0+708] <= intermediate[4095+708:0+708] + a; end
12'd709: begin if(a[709]==1) 
	 		intermediate[4095+709:0+709] <= intermediate[4095+709:0+709] + a; end
12'd710: begin if(a[710]==1) 
	 		intermediate[4095+710:0+710] <= intermediate[4095+710:0+710] + a; end
12'd711: begin if(a[711]==1) 
	 		intermediate[4095+711:0+711] <= intermediate[4095+711:0+711] + a; end
12'd712: begin if(a[712]==1) 
	 		intermediate[4095+712:0+712] <= intermediate[4095+712:0+712] + a; end
12'd713: begin if(a[713]==1) 
	 		intermediate[4095+713:0+713] <= intermediate[4095+713:0+713] + a; end
12'd714: begin if(a[714]==1) 
	 		intermediate[4095+714:0+714] <= intermediate[4095+714:0+714] + a; end
12'd715: begin if(a[715]==1) 
	 		intermediate[4095+715:0+715] <= intermediate[4095+715:0+715] + a; end
12'd716: begin if(a[716]==1) 
	 		intermediate[4095+716:0+716] <= intermediate[4095+716:0+716] + a; end
12'd717: begin if(a[717]==1) 
	 		intermediate[4095+717:0+717] <= intermediate[4095+717:0+717] + a; end
12'd718: begin if(a[718]==1) 
	 		intermediate[4095+718:0+718] <= intermediate[4095+718:0+718] + a; end
12'd719: begin if(a[719]==1) 
	 		intermediate[4095+719:0+719] <= intermediate[4095+719:0+719] + a; end
12'd720: begin if(a[720]==1) 
	 		intermediate[4095+720:0+720] <= intermediate[4095+720:0+720] + a; end
12'd721: begin if(a[721]==1) 
	 		intermediate[4095+721:0+721] <= intermediate[4095+721:0+721] + a; end
12'd722: begin if(a[722]==1) 
	 		intermediate[4095+722:0+722] <= intermediate[4095+722:0+722] + a; end
12'd723: begin if(a[723]==1) 
	 		intermediate[4095+723:0+723] <= intermediate[4095+723:0+723] + a; end
12'd724: begin if(a[724]==1) 
	 		intermediate[4095+724:0+724] <= intermediate[4095+724:0+724] + a; end
12'd725: begin if(a[725]==1) 
	 		intermediate[4095+725:0+725] <= intermediate[4095+725:0+725] + a; end
12'd726: begin if(a[726]==1) 
	 		intermediate[4095+726:0+726] <= intermediate[4095+726:0+726] + a; end
12'd727: begin if(a[727]==1) 
	 		intermediate[4095+727:0+727] <= intermediate[4095+727:0+727] + a; end
12'd728: begin if(a[728]==1) 
	 		intermediate[4095+728:0+728] <= intermediate[4095+728:0+728] + a; end
12'd729: begin if(a[729]==1) 
	 		intermediate[4095+729:0+729] <= intermediate[4095+729:0+729] + a; end
12'd730: begin if(a[730]==1) 
	 		intermediate[4095+730:0+730] <= intermediate[4095+730:0+730] + a; end
12'd731: begin if(a[731]==1) 
	 		intermediate[4095+731:0+731] <= intermediate[4095+731:0+731] + a; end
12'd732: begin if(a[732]==1) 
	 		intermediate[4095+732:0+732] <= intermediate[4095+732:0+732] + a; end
12'd733: begin if(a[733]==1) 
	 		intermediate[4095+733:0+733] <= intermediate[4095+733:0+733] + a; end
12'd734: begin if(a[734]==1) 
	 		intermediate[4095+734:0+734] <= intermediate[4095+734:0+734] + a; end
12'd735: begin if(a[735]==1) 
	 		intermediate[4095+735:0+735] <= intermediate[4095+735:0+735] + a; end
12'd736: begin if(a[736]==1) 
	 		intermediate[4095+736:0+736] <= intermediate[4095+736:0+736] + a; end
12'd737: begin if(a[737]==1) 
	 		intermediate[4095+737:0+737] <= intermediate[4095+737:0+737] + a; end
12'd738: begin if(a[738]==1) 
	 		intermediate[4095+738:0+738] <= intermediate[4095+738:0+738] + a; end
12'd739: begin if(a[739]==1) 
	 		intermediate[4095+739:0+739] <= intermediate[4095+739:0+739] + a; end
12'd740: begin if(a[740]==1) 
	 		intermediate[4095+740:0+740] <= intermediate[4095+740:0+740] + a; end
12'd741: begin if(a[741]==1) 
	 		intermediate[4095+741:0+741] <= intermediate[4095+741:0+741] + a; end
12'd742: begin if(a[742]==1) 
	 		intermediate[4095+742:0+742] <= intermediate[4095+742:0+742] + a; end
12'd743: begin if(a[743]==1) 
	 		intermediate[4095+743:0+743] <= intermediate[4095+743:0+743] + a; end
12'd744: begin if(a[744]==1) 
	 		intermediate[4095+744:0+744] <= intermediate[4095+744:0+744] + a; end
12'd745: begin if(a[745]==1) 
	 		intermediate[4095+745:0+745] <= intermediate[4095+745:0+745] + a; end
12'd746: begin if(a[746]==1) 
	 		intermediate[4095+746:0+746] <= intermediate[4095+746:0+746] + a; end
12'd747: begin if(a[747]==1) 
	 		intermediate[4095+747:0+747] <= intermediate[4095+747:0+747] + a; end
12'd748: begin if(a[748]==1) 
	 		intermediate[4095+748:0+748] <= intermediate[4095+748:0+748] + a; end
12'd749: begin if(a[749]==1) 
	 		intermediate[4095+749:0+749] <= intermediate[4095+749:0+749] + a; end
12'd750: begin if(a[750]==1) 
	 		intermediate[4095+750:0+750] <= intermediate[4095+750:0+750] + a; end
12'd751: begin if(a[751]==1) 
	 		intermediate[4095+751:0+751] <= intermediate[4095+751:0+751] + a; end
12'd752: begin if(a[752]==1) 
	 		intermediate[4095+752:0+752] <= intermediate[4095+752:0+752] + a; end
12'd753: begin if(a[753]==1) 
	 		intermediate[4095+753:0+753] <= intermediate[4095+753:0+753] + a; end
12'd754: begin if(a[754]==1) 
	 		intermediate[4095+754:0+754] <= intermediate[4095+754:0+754] + a; end
12'd755: begin if(a[755]==1) 
	 		intermediate[4095+755:0+755] <= intermediate[4095+755:0+755] + a; end
12'd756: begin if(a[756]==1) 
	 		intermediate[4095+756:0+756] <= intermediate[4095+756:0+756] + a; end
12'd757: begin if(a[757]==1) 
	 		intermediate[4095+757:0+757] <= intermediate[4095+757:0+757] + a; end
12'd758: begin if(a[758]==1) 
	 		intermediate[4095+758:0+758] <= intermediate[4095+758:0+758] + a; end
12'd759: begin if(a[759]==1) 
	 		intermediate[4095+759:0+759] <= intermediate[4095+759:0+759] + a; end
12'd760: begin if(a[760]==1) 
	 		intermediate[4095+760:0+760] <= intermediate[4095+760:0+760] + a; end
12'd761: begin if(a[761]==1) 
	 		intermediate[4095+761:0+761] <= intermediate[4095+761:0+761] + a; end
12'd762: begin if(a[762]==1) 
	 		intermediate[4095+762:0+762] <= intermediate[4095+762:0+762] + a; end
12'd763: begin if(a[763]==1) 
	 		intermediate[4095+763:0+763] <= intermediate[4095+763:0+763] + a; end
12'd764: begin if(a[764]==1) 
	 		intermediate[4095+764:0+764] <= intermediate[4095+764:0+764] + a; end
12'd765: begin if(a[765]==1) 
	 		intermediate[4095+765:0+765] <= intermediate[4095+765:0+765] + a; end
12'd766: begin if(a[766]==1) 
	 		intermediate[4095+766:0+766] <= intermediate[4095+766:0+766] + a; end
12'd767: begin if(a[767]==1) 
	 		intermediate[4095+767:0+767] <= intermediate[4095+767:0+767] + a; end
12'd768: begin if(a[768]==1) 
	 		intermediate[4095+768:0+768] <= intermediate[4095+768:0+768] + a; end
12'd769: begin if(a[769]==1) 
	 		intermediate[4095+769:0+769] <= intermediate[4095+769:0+769] + a; end
12'd770: begin if(a[770]==1) 
	 		intermediate[4095+770:0+770] <= intermediate[4095+770:0+770] + a; end
12'd771: begin if(a[771]==1) 
	 		intermediate[4095+771:0+771] <= intermediate[4095+771:0+771] + a; end
12'd772: begin if(a[772]==1) 
	 		intermediate[4095+772:0+772] <= intermediate[4095+772:0+772] + a; end
12'd773: begin if(a[773]==1) 
	 		intermediate[4095+773:0+773] <= intermediate[4095+773:0+773] + a; end
12'd774: begin if(a[774]==1) 
	 		intermediate[4095+774:0+774] <= intermediate[4095+774:0+774] + a; end
12'd775: begin if(a[775]==1) 
	 		intermediate[4095+775:0+775] <= intermediate[4095+775:0+775] + a; end
12'd776: begin if(a[776]==1) 
	 		intermediate[4095+776:0+776] <= intermediate[4095+776:0+776] + a; end
12'd777: begin if(a[777]==1) 
	 		intermediate[4095+777:0+777] <= intermediate[4095+777:0+777] + a; end
12'd778: begin if(a[778]==1) 
	 		intermediate[4095+778:0+778] <= intermediate[4095+778:0+778] + a; end
12'd779: begin if(a[779]==1) 
	 		intermediate[4095+779:0+779] <= intermediate[4095+779:0+779] + a; end
12'd780: begin if(a[780]==1) 
	 		intermediate[4095+780:0+780] <= intermediate[4095+780:0+780] + a; end
12'd781: begin if(a[781]==1) 
	 		intermediate[4095+781:0+781] <= intermediate[4095+781:0+781] + a; end
12'd782: begin if(a[782]==1) 
	 		intermediate[4095+782:0+782] <= intermediate[4095+782:0+782] + a; end
12'd783: begin if(a[783]==1) 
	 		intermediate[4095+783:0+783] <= intermediate[4095+783:0+783] + a; end
12'd784: begin if(a[784]==1) 
	 		intermediate[4095+784:0+784] <= intermediate[4095+784:0+784] + a; end
12'd785: begin if(a[785]==1) 
	 		intermediate[4095+785:0+785] <= intermediate[4095+785:0+785] + a; end
12'd786: begin if(a[786]==1) 
	 		intermediate[4095+786:0+786] <= intermediate[4095+786:0+786] + a; end
12'd787: begin if(a[787]==1) 
	 		intermediate[4095+787:0+787] <= intermediate[4095+787:0+787] + a; end
12'd788: begin if(a[788]==1) 
	 		intermediate[4095+788:0+788] <= intermediate[4095+788:0+788] + a; end
12'd789: begin if(a[789]==1) 
	 		intermediate[4095+789:0+789] <= intermediate[4095+789:0+789] + a; end
12'd790: begin if(a[790]==1) 
	 		intermediate[4095+790:0+790] <= intermediate[4095+790:0+790] + a; end
12'd791: begin if(a[791]==1) 
	 		intermediate[4095+791:0+791] <= intermediate[4095+791:0+791] + a; end
12'd792: begin if(a[792]==1) 
	 		intermediate[4095+792:0+792] <= intermediate[4095+792:0+792] + a; end
12'd793: begin if(a[793]==1) 
	 		intermediate[4095+793:0+793] <= intermediate[4095+793:0+793] + a; end
12'd794: begin if(a[794]==1) 
	 		intermediate[4095+794:0+794] <= intermediate[4095+794:0+794] + a; end
12'd795: begin if(a[795]==1) 
	 		intermediate[4095+795:0+795] <= intermediate[4095+795:0+795] + a; end
12'd796: begin if(a[796]==1) 
	 		intermediate[4095+796:0+796] <= intermediate[4095+796:0+796] + a; end
12'd797: begin if(a[797]==1) 
	 		intermediate[4095+797:0+797] <= intermediate[4095+797:0+797] + a; end
12'd798: begin if(a[798]==1) 
	 		intermediate[4095+798:0+798] <= intermediate[4095+798:0+798] + a; end
12'd799: begin if(a[799]==1) 
	 		intermediate[4095+799:0+799] <= intermediate[4095+799:0+799] + a; end
12'd800: begin if(a[800]==1) 
	 		intermediate[4095+800:0+800] <= intermediate[4095+800:0+800] + a; end
12'd801: begin if(a[801]==1) 
	 		intermediate[4095+801:0+801] <= intermediate[4095+801:0+801] + a; end
12'd802: begin if(a[802]==1) 
	 		intermediate[4095+802:0+802] <= intermediate[4095+802:0+802] + a; end
12'd803: begin if(a[803]==1) 
	 		intermediate[4095+803:0+803] <= intermediate[4095+803:0+803] + a; end
12'd804: begin if(a[804]==1) 
	 		intermediate[4095+804:0+804] <= intermediate[4095+804:0+804] + a; end
12'd805: begin if(a[805]==1) 
	 		intermediate[4095+805:0+805] <= intermediate[4095+805:0+805] + a; end
12'd806: begin if(a[806]==1) 
	 		intermediate[4095+806:0+806] <= intermediate[4095+806:0+806] + a; end
12'd807: begin if(a[807]==1) 
	 		intermediate[4095+807:0+807] <= intermediate[4095+807:0+807] + a; end
12'd808: begin if(a[808]==1) 
	 		intermediate[4095+808:0+808] <= intermediate[4095+808:0+808] + a; end
12'd809: begin if(a[809]==1) 
	 		intermediate[4095+809:0+809] <= intermediate[4095+809:0+809] + a; end
12'd810: begin if(a[810]==1) 
	 		intermediate[4095+810:0+810] <= intermediate[4095+810:0+810] + a; end
12'd811: begin if(a[811]==1) 
	 		intermediate[4095+811:0+811] <= intermediate[4095+811:0+811] + a; end
12'd812: begin if(a[812]==1) 
	 		intermediate[4095+812:0+812] <= intermediate[4095+812:0+812] + a; end
12'd813: begin if(a[813]==1) 
	 		intermediate[4095+813:0+813] <= intermediate[4095+813:0+813] + a; end
12'd814: begin if(a[814]==1) 
	 		intermediate[4095+814:0+814] <= intermediate[4095+814:0+814] + a; end
12'd815: begin if(a[815]==1) 
	 		intermediate[4095+815:0+815] <= intermediate[4095+815:0+815] + a; end
12'd816: begin if(a[816]==1) 
	 		intermediate[4095+816:0+816] <= intermediate[4095+816:0+816] + a; end
12'd817: begin if(a[817]==1) 
	 		intermediate[4095+817:0+817] <= intermediate[4095+817:0+817] + a; end
12'd818: begin if(a[818]==1) 
	 		intermediate[4095+818:0+818] <= intermediate[4095+818:0+818] + a; end
12'd819: begin if(a[819]==1) 
	 		intermediate[4095+819:0+819] <= intermediate[4095+819:0+819] + a; end
12'd820: begin if(a[820]==1) 
	 		intermediate[4095+820:0+820] <= intermediate[4095+820:0+820] + a; end
12'd821: begin if(a[821]==1) 
	 		intermediate[4095+821:0+821] <= intermediate[4095+821:0+821] + a; end
12'd822: begin if(a[822]==1) 
	 		intermediate[4095+822:0+822] <= intermediate[4095+822:0+822] + a; end
12'd823: begin if(a[823]==1) 
	 		intermediate[4095+823:0+823] <= intermediate[4095+823:0+823] + a; end
12'd824: begin if(a[824]==1) 
	 		intermediate[4095+824:0+824] <= intermediate[4095+824:0+824] + a; end
12'd825: begin if(a[825]==1) 
	 		intermediate[4095+825:0+825] <= intermediate[4095+825:0+825] + a; end
12'd826: begin if(a[826]==1) 
	 		intermediate[4095+826:0+826] <= intermediate[4095+826:0+826] + a; end
12'd827: begin if(a[827]==1) 
	 		intermediate[4095+827:0+827] <= intermediate[4095+827:0+827] + a; end
12'd828: begin if(a[828]==1) 
	 		intermediate[4095+828:0+828] <= intermediate[4095+828:0+828] + a; end
12'd829: begin if(a[829]==1) 
	 		intermediate[4095+829:0+829] <= intermediate[4095+829:0+829] + a; end
12'd830: begin if(a[830]==1) 
	 		intermediate[4095+830:0+830] <= intermediate[4095+830:0+830] + a; end
12'd831: begin if(a[831]==1) 
	 		intermediate[4095+831:0+831] <= intermediate[4095+831:0+831] + a; end
12'd832: begin if(a[832]==1) 
	 		intermediate[4095+832:0+832] <= intermediate[4095+832:0+832] + a; end
12'd833: begin if(a[833]==1) 
	 		intermediate[4095+833:0+833] <= intermediate[4095+833:0+833] + a; end
12'd834: begin if(a[834]==1) 
	 		intermediate[4095+834:0+834] <= intermediate[4095+834:0+834] + a; end
12'd835: begin if(a[835]==1) 
	 		intermediate[4095+835:0+835] <= intermediate[4095+835:0+835] + a; end
12'd836: begin if(a[836]==1) 
	 		intermediate[4095+836:0+836] <= intermediate[4095+836:0+836] + a; end
12'd837: begin if(a[837]==1) 
	 		intermediate[4095+837:0+837] <= intermediate[4095+837:0+837] + a; end
12'd838: begin if(a[838]==1) 
	 		intermediate[4095+838:0+838] <= intermediate[4095+838:0+838] + a; end
12'd839: begin if(a[839]==1) 
	 		intermediate[4095+839:0+839] <= intermediate[4095+839:0+839] + a; end
12'd840: begin if(a[840]==1) 
	 		intermediate[4095+840:0+840] <= intermediate[4095+840:0+840] + a; end
12'd841: begin if(a[841]==1) 
	 		intermediate[4095+841:0+841] <= intermediate[4095+841:0+841] + a; end
12'd842: begin if(a[842]==1) 
	 		intermediate[4095+842:0+842] <= intermediate[4095+842:0+842] + a; end
12'd843: begin if(a[843]==1) 
	 		intermediate[4095+843:0+843] <= intermediate[4095+843:0+843] + a; end
12'd844: begin if(a[844]==1) 
	 		intermediate[4095+844:0+844] <= intermediate[4095+844:0+844] + a; end
12'd845: begin if(a[845]==1) 
	 		intermediate[4095+845:0+845] <= intermediate[4095+845:0+845] + a; end
12'd846: begin if(a[846]==1) 
	 		intermediate[4095+846:0+846] <= intermediate[4095+846:0+846] + a; end
12'd847: begin if(a[847]==1) 
	 		intermediate[4095+847:0+847] <= intermediate[4095+847:0+847] + a; end
12'd848: begin if(a[848]==1) 
	 		intermediate[4095+848:0+848] <= intermediate[4095+848:0+848] + a; end
12'd849: begin if(a[849]==1) 
	 		intermediate[4095+849:0+849] <= intermediate[4095+849:0+849] + a; end
12'd850: begin if(a[850]==1) 
	 		intermediate[4095+850:0+850] <= intermediate[4095+850:0+850] + a; end
12'd851: begin if(a[851]==1) 
	 		intermediate[4095+851:0+851] <= intermediate[4095+851:0+851] + a; end
12'd852: begin if(a[852]==1) 
	 		intermediate[4095+852:0+852] <= intermediate[4095+852:0+852] + a; end
12'd853: begin if(a[853]==1) 
	 		intermediate[4095+853:0+853] <= intermediate[4095+853:0+853] + a; end
12'd854: begin if(a[854]==1) 
	 		intermediate[4095+854:0+854] <= intermediate[4095+854:0+854] + a; end
12'd855: begin if(a[855]==1) 
	 		intermediate[4095+855:0+855] <= intermediate[4095+855:0+855] + a; end
12'd856: begin if(a[856]==1) 
	 		intermediate[4095+856:0+856] <= intermediate[4095+856:0+856] + a; end
12'd857: begin if(a[857]==1) 
	 		intermediate[4095+857:0+857] <= intermediate[4095+857:0+857] + a; end
12'd858: begin if(a[858]==1) 
	 		intermediate[4095+858:0+858] <= intermediate[4095+858:0+858] + a; end
12'd859: begin if(a[859]==1) 
	 		intermediate[4095+859:0+859] <= intermediate[4095+859:0+859] + a; end
12'd860: begin if(a[860]==1) 
	 		intermediate[4095+860:0+860] <= intermediate[4095+860:0+860] + a; end
12'd861: begin if(a[861]==1) 
	 		intermediate[4095+861:0+861] <= intermediate[4095+861:0+861] + a; end
12'd862: begin if(a[862]==1) 
	 		intermediate[4095+862:0+862] <= intermediate[4095+862:0+862] + a; end
12'd863: begin if(a[863]==1) 
	 		intermediate[4095+863:0+863] <= intermediate[4095+863:0+863] + a; end
12'd864: begin if(a[864]==1) 
	 		intermediate[4095+864:0+864] <= intermediate[4095+864:0+864] + a; end
12'd865: begin if(a[865]==1) 
	 		intermediate[4095+865:0+865] <= intermediate[4095+865:0+865] + a; end
12'd866: begin if(a[866]==1) 
	 		intermediate[4095+866:0+866] <= intermediate[4095+866:0+866] + a; end
12'd867: begin if(a[867]==1) 
	 		intermediate[4095+867:0+867] <= intermediate[4095+867:0+867] + a; end
12'd868: begin if(a[868]==1) 
	 		intermediate[4095+868:0+868] <= intermediate[4095+868:0+868] + a; end
12'd869: begin if(a[869]==1) 
	 		intermediate[4095+869:0+869] <= intermediate[4095+869:0+869] + a; end
12'd870: begin if(a[870]==1) 
	 		intermediate[4095+870:0+870] <= intermediate[4095+870:0+870] + a; end
12'd871: begin if(a[871]==1) 
	 		intermediate[4095+871:0+871] <= intermediate[4095+871:0+871] + a; end
12'd872: begin if(a[872]==1) 
	 		intermediate[4095+872:0+872] <= intermediate[4095+872:0+872] + a; end
12'd873: begin if(a[873]==1) 
	 		intermediate[4095+873:0+873] <= intermediate[4095+873:0+873] + a; end
12'd874: begin if(a[874]==1) 
	 		intermediate[4095+874:0+874] <= intermediate[4095+874:0+874] + a; end
12'd875: begin if(a[875]==1) 
	 		intermediate[4095+875:0+875] <= intermediate[4095+875:0+875] + a; end
12'd876: begin if(a[876]==1) 
	 		intermediate[4095+876:0+876] <= intermediate[4095+876:0+876] + a; end
12'd877: begin if(a[877]==1) 
	 		intermediate[4095+877:0+877] <= intermediate[4095+877:0+877] + a; end
12'd878: begin if(a[878]==1) 
	 		intermediate[4095+878:0+878] <= intermediate[4095+878:0+878] + a; end
12'd879: begin if(a[879]==1) 
	 		intermediate[4095+879:0+879] <= intermediate[4095+879:0+879] + a; end
12'd880: begin if(a[880]==1) 
	 		intermediate[4095+880:0+880] <= intermediate[4095+880:0+880] + a; end
12'd881: begin if(a[881]==1) 
	 		intermediate[4095+881:0+881] <= intermediate[4095+881:0+881] + a; end
12'd882: begin if(a[882]==1) 
	 		intermediate[4095+882:0+882] <= intermediate[4095+882:0+882] + a; end
12'd883: begin if(a[883]==1) 
	 		intermediate[4095+883:0+883] <= intermediate[4095+883:0+883] + a; end
12'd884: begin if(a[884]==1) 
	 		intermediate[4095+884:0+884] <= intermediate[4095+884:0+884] + a; end
12'd885: begin if(a[885]==1) 
	 		intermediate[4095+885:0+885] <= intermediate[4095+885:0+885] + a; end
12'd886: begin if(a[886]==1) 
	 		intermediate[4095+886:0+886] <= intermediate[4095+886:0+886] + a; end
12'd887: begin if(a[887]==1) 
	 		intermediate[4095+887:0+887] <= intermediate[4095+887:0+887] + a; end
12'd888: begin if(a[888]==1) 
	 		intermediate[4095+888:0+888] <= intermediate[4095+888:0+888] + a; end
12'd889: begin if(a[889]==1) 
	 		intermediate[4095+889:0+889] <= intermediate[4095+889:0+889] + a; end
12'd890: begin if(a[890]==1) 
	 		intermediate[4095+890:0+890] <= intermediate[4095+890:0+890] + a; end
12'd891: begin if(a[891]==1) 
	 		intermediate[4095+891:0+891] <= intermediate[4095+891:0+891] + a; end
12'd892: begin if(a[892]==1) 
	 		intermediate[4095+892:0+892] <= intermediate[4095+892:0+892] + a; end
12'd893: begin if(a[893]==1) 
	 		intermediate[4095+893:0+893] <= intermediate[4095+893:0+893] + a; end
12'd894: begin if(a[894]==1) 
	 		intermediate[4095+894:0+894] <= intermediate[4095+894:0+894] + a; end
12'd895: begin if(a[895]==1) 
	 		intermediate[4095+895:0+895] <= intermediate[4095+895:0+895] + a; end
12'd896: begin if(a[896]==1) 
	 		intermediate[4095+896:0+896] <= intermediate[4095+896:0+896] + a; end
12'd897: begin if(a[897]==1) 
	 		intermediate[4095+897:0+897] <= intermediate[4095+897:0+897] + a; end
12'd898: begin if(a[898]==1) 
	 		intermediate[4095+898:0+898] <= intermediate[4095+898:0+898] + a; end
12'd899: begin if(a[899]==1) 
	 		intermediate[4095+899:0+899] <= intermediate[4095+899:0+899] + a; end
12'd900: begin if(a[900]==1) 
	 		intermediate[4095+900:0+900] <= intermediate[4095+900:0+900] + a; end
12'd901: begin if(a[901]==1) 
	 		intermediate[4095+901:0+901] <= intermediate[4095+901:0+901] + a; end
12'd902: begin if(a[902]==1) 
	 		intermediate[4095+902:0+902] <= intermediate[4095+902:0+902] + a; end
12'd903: begin if(a[903]==1) 
	 		intermediate[4095+903:0+903] <= intermediate[4095+903:0+903] + a; end
12'd904: begin if(a[904]==1) 
	 		intermediate[4095+904:0+904] <= intermediate[4095+904:0+904] + a; end
12'd905: begin if(a[905]==1) 
	 		intermediate[4095+905:0+905] <= intermediate[4095+905:0+905] + a; end
12'd906: begin if(a[906]==1) 
	 		intermediate[4095+906:0+906] <= intermediate[4095+906:0+906] + a; end
12'd907: begin if(a[907]==1) 
	 		intermediate[4095+907:0+907] <= intermediate[4095+907:0+907] + a; end
12'd908: begin if(a[908]==1) 
	 		intermediate[4095+908:0+908] <= intermediate[4095+908:0+908] + a; end
12'd909: begin if(a[909]==1) 
	 		intermediate[4095+909:0+909] <= intermediate[4095+909:0+909] + a; end
12'd910: begin if(a[910]==1) 
	 		intermediate[4095+910:0+910] <= intermediate[4095+910:0+910] + a; end
12'd911: begin if(a[911]==1) 
	 		intermediate[4095+911:0+911] <= intermediate[4095+911:0+911] + a; end
12'd912: begin if(a[912]==1) 
	 		intermediate[4095+912:0+912] <= intermediate[4095+912:0+912] + a; end
12'd913: begin if(a[913]==1) 
	 		intermediate[4095+913:0+913] <= intermediate[4095+913:0+913] + a; end
12'd914: begin if(a[914]==1) 
	 		intermediate[4095+914:0+914] <= intermediate[4095+914:0+914] + a; end
12'd915: begin if(a[915]==1) 
	 		intermediate[4095+915:0+915] <= intermediate[4095+915:0+915] + a; end
12'd916: begin if(a[916]==1) 
	 		intermediate[4095+916:0+916] <= intermediate[4095+916:0+916] + a; end
12'd917: begin if(a[917]==1) 
	 		intermediate[4095+917:0+917] <= intermediate[4095+917:0+917] + a; end
12'd918: begin if(a[918]==1) 
	 		intermediate[4095+918:0+918] <= intermediate[4095+918:0+918] + a; end
12'd919: begin if(a[919]==1) 
	 		intermediate[4095+919:0+919] <= intermediate[4095+919:0+919] + a; end
12'd920: begin if(a[920]==1) 
	 		intermediate[4095+920:0+920] <= intermediate[4095+920:0+920] + a; end
12'd921: begin if(a[921]==1) 
	 		intermediate[4095+921:0+921] <= intermediate[4095+921:0+921] + a; end
12'd922: begin if(a[922]==1) 
	 		intermediate[4095+922:0+922] <= intermediate[4095+922:0+922] + a; end
12'd923: begin if(a[923]==1) 
	 		intermediate[4095+923:0+923] <= intermediate[4095+923:0+923] + a; end
12'd924: begin if(a[924]==1) 
	 		intermediate[4095+924:0+924] <= intermediate[4095+924:0+924] + a; end
12'd925: begin if(a[925]==1) 
	 		intermediate[4095+925:0+925] <= intermediate[4095+925:0+925] + a; end
12'd926: begin if(a[926]==1) 
	 		intermediate[4095+926:0+926] <= intermediate[4095+926:0+926] + a; end
12'd927: begin if(a[927]==1) 
	 		intermediate[4095+927:0+927] <= intermediate[4095+927:0+927] + a; end
12'd928: begin if(a[928]==1) 
	 		intermediate[4095+928:0+928] <= intermediate[4095+928:0+928] + a; end
12'd929: begin if(a[929]==1) 
	 		intermediate[4095+929:0+929] <= intermediate[4095+929:0+929] + a; end
12'd930: begin if(a[930]==1) 
	 		intermediate[4095+930:0+930] <= intermediate[4095+930:0+930] + a; end
12'd931: begin if(a[931]==1) 
	 		intermediate[4095+931:0+931] <= intermediate[4095+931:0+931] + a; end
12'd932: begin if(a[932]==1) 
	 		intermediate[4095+932:0+932] <= intermediate[4095+932:0+932] + a; end
12'd933: begin if(a[933]==1) 
	 		intermediate[4095+933:0+933] <= intermediate[4095+933:0+933] + a; end
12'd934: begin if(a[934]==1) 
	 		intermediate[4095+934:0+934] <= intermediate[4095+934:0+934] + a; end
12'd935: begin if(a[935]==1) 
	 		intermediate[4095+935:0+935] <= intermediate[4095+935:0+935] + a; end
12'd936: begin if(a[936]==1) 
	 		intermediate[4095+936:0+936] <= intermediate[4095+936:0+936] + a; end
12'd937: begin if(a[937]==1) 
	 		intermediate[4095+937:0+937] <= intermediate[4095+937:0+937] + a; end
12'd938: begin if(a[938]==1) 
	 		intermediate[4095+938:0+938] <= intermediate[4095+938:0+938] + a; end
12'd939: begin if(a[939]==1) 
	 		intermediate[4095+939:0+939] <= intermediate[4095+939:0+939] + a; end
12'd940: begin if(a[940]==1) 
	 		intermediate[4095+940:0+940] <= intermediate[4095+940:0+940] + a; end
12'd941: begin if(a[941]==1) 
	 		intermediate[4095+941:0+941] <= intermediate[4095+941:0+941] + a; end
12'd942: begin if(a[942]==1) 
	 		intermediate[4095+942:0+942] <= intermediate[4095+942:0+942] + a; end
12'd943: begin if(a[943]==1) 
	 		intermediate[4095+943:0+943] <= intermediate[4095+943:0+943] + a; end
12'd944: begin if(a[944]==1) 
	 		intermediate[4095+944:0+944] <= intermediate[4095+944:0+944] + a; end
12'd945: begin if(a[945]==1) 
	 		intermediate[4095+945:0+945] <= intermediate[4095+945:0+945] + a; end
12'd946: begin if(a[946]==1) 
	 		intermediate[4095+946:0+946] <= intermediate[4095+946:0+946] + a; end
12'd947: begin if(a[947]==1) 
	 		intermediate[4095+947:0+947] <= intermediate[4095+947:0+947] + a; end
12'd948: begin if(a[948]==1) 
	 		intermediate[4095+948:0+948] <= intermediate[4095+948:0+948] + a; end
12'd949: begin if(a[949]==1) 
	 		intermediate[4095+949:0+949] <= intermediate[4095+949:0+949] + a; end
12'd950: begin if(a[950]==1) 
	 		intermediate[4095+950:0+950] <= intermediate[4095+950:0+950] + a; end
12'd951: begin if(a[951]==1) 
	 		intermediate[4095+951:0+951] <= intermediate[4095+951:0+951] + a; end
12'd952: begin if(a[952]==1) 
	 		intermediate[4095+952:0+952] <= intermediate[4095+952:0+952] + a; end
12'd953: begin if(a[953]==1) 
	 		intermediate[4095+953:0+953] <= intermediate[4095+953:0+953] + a; end
12'd954: begin if(a[954]==1) 
	 		intermediate[4095+954:0+954] <= intermediate[4095+954:0+954] + a; end
12'd955: begin if(a[955]==1) 
	 		intermediate[4095+955:0+955] <= intermediate[4095+955:0+955] + a; end
12'd956: begin if(a[956]==1) 
	 		intermediate[4095+956:0+956] <= intermediate[4095+956:0+956] + a; end
12'd957: begin if(a[957]==1) 
	 		intermediate[4095+957:0+957] <= intermediate[4095+957:0+957] + a; end
12'd958: begin if(a[958]==1) 
	 		intermediate[4095+958:0+958] <= intermediate[4095+958:0+958] + a; end
12'd959: begin if(a[959]==1) 
	 		intermediate[4095+959:0+959] <= intermediate[4095+959:0+959] + a; end
12'd960: begin if(a[960]==1) 
	 		intermediate[4095+960:0+960] <= intermediate[4095+960:0+960] + a; end
12'd961: begin if(a[961]==1) 
	 		intermediate[4095+961:0+961] <= intermediate[4095+961:0+961] + a; end
12'd962: begin if(a[962]==1) 
	 		intermediate[4095+962:0+962] <= intermediate[4095+962:0+962] + a; end
12'd963: begin if(a[963]==1) 
	 		intermediate[4095+963:0+963] <= intermediate[4095+963:0+963] + a; end
12'd964: begin if(a[964]==1) 
	 		intermediate[4095+964:0+964] <= intermediate[4095+964:0+964] + a; end
12'd965: begin if(a[965]==1) 
	 		intermediate[4095+965:0+965] <= intermediate[4095+965:0+965] + a; end
12'd966: begin if(a[966]==1) 
	 		intermediate[4095+966:0+966] <= intermediate[4095+966:0+966] + a; end
12'd967: begin if(a[967]==1) 
	 		intermediate[4095+967:0+967] <= intermediate[4095+967:0+967] + a; end
12'd968: begin if(a[968]==1) 
	 		intermediate[4095+968:0+968] <= intermediate[4095+968:0+968] + a; end
12'd969: begin if(a[969]==1) 
	 		intermediate[4095+969:0+969] <= intermediate[4095+969:0+969] + a; end
12'd970: begin if(a[970]==1) 
	 		intermediate[4095+970:0+970] <= intermediate[4095+970:0+970] + a; end
12'd971: begin if(a[971]==1) 
	 		intermediate[4095+971:0+971] <= intermediate[4095+971:0+971] + a; end
12'd972: begin if(a[972]==1) 
	 		intermediate[4095+972:0+972] <= intermediate[4095+972:0+972] + a; end
12'd973: begin if(a[973]==1) 
	 		intermediate[4095+973:0+973] <= intermediate[4095+973:0+973] + a; end
12'd974: begin if(a[974]==1) 
	 		intermediate[4095+974:0+974] <= intermediate[4095+974:0+974] + a; end
12'd975: begin if(a[975]==1) 
	 		intermediate[4095+975:0+975] <= intermediate[4095+975:0+975] + a; end
12'd976: begin if(a[976]==1) 
	 		intermediate[4095+976:0+976] <= intermediate[4095+976:0+976] + a; end
12'd977: begin if(a[977]==1) 
	 		intermediate[4095+977:0+977] <= intermediate[4095+977:0+977] + a; end
12'd978: begin if(a[978]==1) 
	 		intermediate[4095+978:0+978] <= intermediate[4095+978:0+978] + a; end
12'd979: begin if(a[979]==1) 
	 		intermediate[4095+979:0+979] <= intermediate[4095+979:0+979] + a; end
12'd980: begin if(a[980]==1) 
	 		intermediate[4095+980:0+980] <= intermediate[4095+980:0+980] + a; end
12'd981: begin if(a[981]==1) 
	 		intermediate[4095+981:0+981] <= intermediate[4095+981:0+981] + a; end
12'd982: begin if(a[982]==1) 
	 		intermediate[4095+982:0+982] <= intermediate[4095+982:0+982] + a; end
12'd983: begin if(a[983]==1) 
	 		intermediate[4095+983:0+983] <= intermediate[4095+983:0+983] + a; end
12'd984: begin if(a[984]==1) 
	 		intermediate[4095+984:0+984] <= intermediate[4095+984:0+984] + a; end
12'd985: begin if(a[985]==1) 
	 		intermediate[4095+985:0+985] <= intermediate[4095+985:0+985] + a; end
12'd986: begin if(a[986]==1) 
	 		intermediate[4095+986:0+986] <= intermediate[4095+986:0+986] + a; end
12'd987: begin if(a[987]==1) 
	 		intermediate[4095+987:0+987] <= intermediate[4095+987:0+987] + a; end
12'd988: begin if(a[988]==1) 
	 		intermediate[4095+988:0+988] <= intermediate[4095+988:0+988] + a; end
12'd989: begin if(a[989]==1) 
	 		intermediate[4095+989:0+989] <= intermediate[4095+989:0+989] + a; end
12'd990: begin if(a[990]==1) 
	 		intermediate[4095+990:0+990] <= intermediate[4095+990:0+990] + a; end
12'd991: begin if(a[991]==1) 
	 		intermediate[4095+991:0+991] <= intermediate[4095+991:0+991] + a; end
12'd992: begin if(a[992]==1) 
	 		intermediate[4095+992:0+992] <= intermediate[4095+992:0+992] + a; end
12'd993: begin if(a[993]==1) 
	 		intermediate[4095+993:0+993] <= intermediate[4095+993:0+993] + a; end
12'd994: begin if(a[994]==1) 
	 		intermediate[4095+994:0+994] <= intermediate[4095+994:0+994] + a; end
12'd995: begin if(a[995]==1) 
	 		intermediate[4095+995:0+995] <= intermediate[4095+995:0+995] + a; end
12'd996: begin if(a[996]==1) 
	 		intermediate[4095+996:0+996] <= intermediate[4095+996:0+996] + a; end
12'd997: begin if(a[997]==1) 
	 		intermediate[4095+997:0+997] <= intermediate[4095+997:0+997] + a; end
12'd998: begin if(a[998]==1) 
	 		intermediate[4095+998:0+998] <= intermediate[4095+998:0+998] + a; end
12'd999: begin if(a[999]==1) 
	 		intermediate[4095+999:0+999] <= intermediate[4095+999:0+999] + a; end
12'd1000: begin if(a[1000]==1) 
	 		intermediate[4095+1000:0+1000] <= intermediate[4095+1000:0+1000] + a; end
12'd1001: begin if(a[1001]==1) 
	 		intermediate[4095+1001:0+1001] <= intermediate[4095+1001:0+1001] + a; end
12'd1002: begin if(a[1002]==1) 
	 		intermediate[4095+1002:0+1002] <= intermediate[4095+1002:0+1002] + a; end
12'd1003: begin if(a[1003]==1) 
	 		intermediate[4095+1003:0+1003] <= intermediate[4095+1003:0+1003] + a; end
12'd1004: begin if(a[1004]==1) 
	 		intermediate[4095+1004:0+1004] <= intermediate[4095+1004:0+1004] + a; end
12'd1005: begin if(a[1005]==1) 
	 		intermediate[4095+1005:0+1005] <= intermediate[4095+1005:0+1005] + a; end
12'd1006: begin if(a[1006]==1) 
	 		intermediate[4095+1006:0+1006] <= intermediate[4095+1006:0+1006] + a; end
12'd1007: begin if(a[1007]==1) 
	 		intermediate[4095+1007:0+1007] <= intermediate[4095+1007:0+1007] + a; end
12'd1008: begin if(a[1008]==1) 
	 		intermediate[4095+1008:0+1008] <= intermediate[4095+1008:0+1008] + a; end
12'd1009: begin if(a[1009]==1) 
	 		intermediate[4095+1009:0+1009] <= intermediate[4095+1009:0+1009] + a; end
12'd1010: begin if(a[1010]==1) 
	 		intermediate[4095+1010:0+1010] <= intermediate[4095+1010:0+1010] + a; end
12'd1011: begin if(a[1011]==1) 
	 		intermediate[4095+1011:0+1011] <= intermediate[4095+1011:0+1011] + a; end
12'd1012: begin if(a[1012]==1) 
	 		intermediate[4095+1012:0+1012] <= intermediate[4095+1012:0+1012] + a; end
12'd1013: begin if(a[1013]==1) 
	 		intermediate[4095+1013:0+1013] <= intermediate[4095+1013:0+1013] + a; end
12'd1014: begin if(a[1014]==1) 
	 		intermediate[4095+1014:0+1014] <= intermediate[4095+1014:0+1014] + a; end
12'd1015: begin if(a[1015]==1) 
	 		intermediate[4095+1015:0+1015] <= intermediate[4095+1015:0+1015] + a; end
12'd1016: begin if(a[1016]==1) 
	 		intermediate[4095+1016:0+1016] <= intermediate[4095+1016:0+1016] + a; end
12'd1017: begin if(a[1017]==1) 
	 		intermediate[4095+1017:0+1017] <= intermediate[4095+1017:0+1017] + a; end
12'd1018: begin if(a[1018]==1) 
	 		intermediate[4095+1018:0+1018] <= intermediate[4095+1018:0+1018] + a; end
12'd1019: begin if(a[1019]==1) 
	 		intermediate[4095+1019:0+1019] <= intermediate[4095+1019:0+1019] + a; end
12'd1020: begin if(a[1020]==1) 
	 		intermediate[4095+1020:0+1020] <= intermediate[4095+1020:0+1020] + a; end
12'd1021: begin if(a[1021]==1) 
	 		intermediate[4095+1021:0+1021] <= intermediate[4095+1021:0+1021] + a; end
12'd1022: begin if(a[1022]==1) 
	 		intermediate[4095+1022:0+1022] <= intermediate[4095+1022:0+1022] + a; end
12'd1023: begin if(a[1023]==1) 
	 		intermediate[4095+1023:0+1023] <= intermediate[4095+1023:0+1023] + a; end
12'd1024: begin if(a[1024]==1) 
	 		intermediate[4095+1024:0+1024] <= intermediate[4095+1024:0+1024] + a; end
12'd1025: begin if(a[1025]==1) 
	 		intermediate[4095+1025:0+1025] <= intermediate[4095+1025:0+1025] + a; end
12'd1026: begin if(a[1026]==1) 
	 		intermediate[4095+1026:0+1026] <= intermediate[4095+1026:0+1026] + a; end
12'd1027: begin if(a[1027]==1) 
	 		intermediate[4095+1027:0+1027] <= intermediate[4095+1027:0+1027] + a; end
12'd1028: begin if(a[1028]==1) 
	 		intermediate[4095+1028:0+1028] <= intermediate[4095+1028:0+1028] + a; end
12'd1029: begin if(a[1029]==1) 
	 		intermediate[4095+1029:0+1029] <= intermediate[4095+1029:0+1029] + a; end
12'd1030: begin if(a[1030]==1) 
	 		intermediate[4095+1030:0+1030] <= intermediate[4095+1030:0+1030] + a; end
12'd1031: begin if(a[1031]==1) 
	 		intermediate[4095+1031:0+1031] <= intermediate[4095+1031:0+1031] + a; end
12'd1032: begin if(a[1032]==1) 
	 		intermediate[4095+1032:0+1032] <= intermediate[4095+1032:0+1032] + a; end
12'd1033: begin if(a[1033]==1) 
	 		intermediate[4095+1033:0+1033] <= intermediate[4095+1033:0+1033] + a; end
12'd1034: begin if(a[1034]==1) 
	 		intermediate[4095+1034:0+1034] <= intermediate[4095+1034:0+1034] + a; end
12'd1035: begin if(a[1035]==1) 
	 		intermediate[4095+1035:0+1035] <= intermediate[4095+1035:0+1035] + a; end
12'd1036: begin if(a[1036]==1) 
	 		intermediate[4095+1036:0+1036] <= intermediate[4095+1036:0+1036] + a; end
12'd1037: begin if(a[1037]==1) 
	 		intermediate[4095+1037:0+1037] <= intermediate[4095+1037:0+1037] + a; end
12'd1038: begin if(a[1038]==1) 
	 		intermediate[4095+1038:0+1038] <= intermediate[4095+1038:0+1038] + a; end
12'd1039: begin if(a[1039]==1) 
	 		intermediate[4095+1039:0+1039] <= intermediate[4095+1039:0+1039] + a; end
12'd1040: begin if(a[1040]==1) 
	 		intermediate[4095+1040:0+1040] <= intermediate[4095+1040:0+1040] + a; end
12'd1041: begin if(a[1041]==1) 
	 		intermediate[4095+1041:0+1041] <= intermediate[4095+1041:0+1041] + a; end
12'd1042: begin if(a[1042]==1) 
	 		intermediate[4095+1042:0+1042] <= intermediate[4095+1042:0+1042] + a; end
12'd1043: begin if(a[1043]==1) 
	 		intermediate[4095+1043:0+1043] <= intermediate[4095+1043:0+1043] + a; end
12'd1044: begin if(a[1044]==1) 
	 		intermediate[4095+1044:0+1044] <= intermediate[4095+1044:0+1044] + a; end
12'd1045: begin if(a[1045]==1) 
	 		intermediate[4095+1045:0+1045] <= intermediate[4095+1045:0+1045] + a; end
12'd1046: begin if(a[1046]==1) 
	 		intermediate[4095+1046:0+1046] <= intermediate[4095+1046:0+1046] + a; end
12'd1047: begin if(a[1047]==1) 
	 		intermediate[4095+1047:0+1047] <= intermediate[4095+1047:0+1047] + a; end
12'd1048: begin if(a[1048]==1) 
	 		intermediate[4095+1048:0+1048] <= intermediate[4095+1048:0+1048] + a; end
12'd1049: begin if(a[1049]==1) 
	 		intermediate[4095+1049:0+1049] <= intermediate[4095+1049:0+1049] + a; end
12'd1050: begin if(a[1050]==1) 
	 		intermediate[4095+1050:0+1050] <= intermediate[4095+1050:0+1050] + a; end
12'd1051: begin if(a[1051]==1) 
	 		intermediate[4095+1051:0+1051] <= intermediate[4095+1051:0+1051] + a; end
12'd1052: begin if(a[1052]==1) 
	 		intermediate[4095+1052:0+1052] <= intermediate[4095+1052:0+1052] + a; end
12'd1053: begin if(a[1053]==1) 
	 		intermediate[4095+1053:0+1053] <= intermediate[4095+1053:0+1053] + a; end
12'd1054: begin if(a[1054]==1) 
	 		intermediate[4095+1054:0+1054] <= intermediate[4095+1054:0+1054] + a; end
12'd1055: begin if(a[1055]==1) 
	 		intermediate[4095+1055:0+1055] <= intermediate[4095+1055:0+1055] + a; end
12'd1056: begin if(a[1056]==1) 
	 		intermediate[4095+1056:0+1056] <= intermediate[4095+1056:0+1056] + a; end
12'd1057: begin if(a[1057]==1) 
	 		intermediate[4095+1057:0+1057] <= intermediate[4095+1057:0+1057] + a; end
12'd1058: begin if(a[1058]==1) 
	 		intermediate[4095+1058:0+1058] <= intermediate[4095+1058:0+1058] + a; end
12'd1059: begin if(a[1059]==1) 
	 		intermediate[4095+1059:0+1059] <= intermediate[4095+1059:0+1059] + a; end
12'd1060: begin if(a[1060]==1) 
	 		intermediate[4095+1060:0+1060] <= intermediate[4095+1060:0+1060] + a; end
12'd1061: begin if(a[1061]==1) 
	 		intermediate[4095+1061:0+1061] <= intermediate[4095+1061:0+1061] + a; end
12'd1062: begin if(a[1062]==1) 
	 		intermediate[4095+1062:0+1062] <= intermediate[4095+1062:0+1062] + a; end
12'd1063: begin if(a[1063]==1) 
	 		intermediate[4095+1063:0+1063] <= intermediate[4095+1063:0+1063] + a; end
12'd1064: begin if(a[1064]==1) 
	 		intermediate[4095+1064:0+1064] <= intermediate[4095+1064:0+1064] + a; end
12'd1065: begin if(a[1065]==1) 
	 		intermediate[4095+1065:0+1065] <= intermediate[4095+1065:0+1065] + a; end
12'd1066: begin if(a[1066]==1) 
	 		intermediate[4095+1066:0+1066] <= intermediate[4095+1066:0+1066] + a; end
12'd1067: begin if(a[1067]==1) 
	 		intermediate[4095+1067:0+1067] <= intermediate[4095+1067:0+1067] + a; end
12'd1068: begin if(a[1068]==1) 
	 		intermediate[4095+1068:0+1068] <= intermediate[4095+1068:0+1068] + a; end
12'd1069: begin if(a[1069]==1) 
	 		intermediate[4095+1069:0+1069] <= intermediate[4095+1069:0+1069] + a; end
12'd1070: begin if(a[1070]==1) 
	 		intermediate[4095+1070:0+1070] <= intermediate[4095+1070:0+1070] + a; end
12'd1071: begin if(a[1071]==1) 
	 		intermediate[4095+1071:0+1071] <= intermediate[4095+1071:0+1071] + a; end
12'd1072: begin if(a[1072]==1) 
	 		intermediate[4095+1072:0+1072] <= intermediate[4095+1072:0+1072] + a; end
12'd1073: begin if(a[1073]==1) 
	 		intermediate[4095+1073:0+1073] <= intermediate[4095+1073:0+1073] + a; end
12'd1074: begin if(a[1074]==1) 
	 		intermediate[4095+1074:0+1074] <= intermediate[4095+1074:0+1074] + a; end
12'd1075: begin if(a[1075]==1) 
	 		intermediate[4095+1075:0+1075] <= intermediate[4095+1075:0+1075] + a; end
12'd1076: begin if(a[1076]==1) 
	 		intermediate[4095+1076:0+1076] <= intermediate[4095+1076:0+1076] + a; end
12'd1077: begin if(a[1077]==1) 
	 		intermediate[4095+1077:0+1077] <= intermediate[4095+1077:0+1077] + a; end
12'd1078: begin if(a[1078]==1) 
	 		intermediate[4095+1078:0+1078] <= intermediate[4095+1078:0+1078] + a; end
12'd1079: begin if(a[1079]==1) 
	 		intermediate[4095+1079:0+1079] <= intermediate[4095+1079:0+1079] + a; end
12'd1080: begin if(a[1080]==1) 
	 		intermediate[4095+1080:0+1080] <= intermediate[4095+1080:0+1080] + a; end
12'd1081: begin if(a[1081]==1) 
	 		intermediate[4095+1081:0+1081] <= intermediate[4095+1081:0+1081] + a; end
12'd1082: begin if(a[1082]==1) 
	 		intermediate[4095+1082:0+1082] <= intermediate[4095+1082:0+1082] + a; end
12'd1083: begin if(a[1083]==1) 
	 		intermediate[4095+1083:0+1083] <= intermediate[4095+1083:0+1083] + a; end
12'd1084: begin if(a[1084]==1) 
	 		intermediate[4095+1084:0+1084] <= intermediate[4095+1084:0+1084] + a; end
12'd1085: begin if(a[1085]==1) 
	 		intermediate[4095+1085:0+1085] <= intermediate[4095+1085:0+1085] + a; end
12'd1086: begin if(a[1086]==1) 
	 		intermediate[4095+1086:0+1086] <= intermediate[4095+1086:0+1086] + a; end
12'd1087: begin if(a[1087]==1) 
	 		intermediate[4095+1087:0+1087] <= intermediate[4095+1087:0+1087] + a; end
12'd1088: begin if(a[1088]==1) 
	 		intermediate[4095+1088:0+1088] <= intermediate[4095+1088:0+1088] + a; end
12'd1089: begin if(a[1089]==1) 
	 		intermediate[4095+1089:0+1089] <= intermediate[4095+1089:0+1089] + a; end
12'd1090: begin if(a[1090]==1) 
	 		intermediate[4095+1090:0+1090] <= intermediate[4095+1090:0+1090] + a; end
12'd1091: begin if(a[1091]==1) 
	 		intermediate[4095+1091:0+1091] <= intermediate[4095+1091:0+1091] + a; end
12'd1092: begin if(a[1092]==1) 
	 		intermediate[4095+1092:0+1092] <= intermediate[4095+1092:0+1092] + a; end
12'd1093: begin if(a[1093]==1) 
	 		intermediate[4095+1093:0+1093] <= intermediate[4095+1093:0+1093] + a; end
12'd1094: begin if(a[1094]==1) 
	 		intermediate[4095+1094:0+1094] <= intermediate[4095+1094:0+1094] + a; end
12'd1095: begin if(a[1095]==1) 
	 		intermediate[4095+1095:0+1095] <= intermediate[4095+1095:0+1095] + a; end
12'd1096: begin if(a[1096]==1) 
	 		intermediate[4095+1096:0+1096] <= intermediate[4095+1096:0+1096] + a; end
12'd1097: begin if(a[1097]==1) 
	 		intermediate[4095+1097:0+1097] <= intermediate[4095+1097:0+1097] + a; end
12'd1098: begin if(a[1098]==1) 
	 		intermediate[4095+1098:0+1098] <= intermediate[4095+1098:0+1098] + a; end
12'd1099: begin if(a[1099]==1) 
	 		intermediate[4095+1099:0+1099] <= intermediate[4095+1099:0+1099] + a; end
12'd1100: begin if(a[1100]==1) 
	 		intermediate[4095+1100:0+1100] <= intermediate[4095+1100:0+1100] + a; end
12'd1101: begin if(a[1101]==1) 
	 		intermediate[4095+1101:0+1101] <= intermediate[4095+1101:0+1101] + a; end
12'd1102: begin if(a[1102]==1) 
	 		intermediate[4095+1102:0+1102] <= intermediate[4095+1102:0+1102] + a; end
12'd1103: begin if(a[1103]==1) 
	 		intermediate[4095+1103:0+1103] <= intermediate[4095+1103:0+1103] + a; end
12'd1104: begin if(a[1104]==1) 
	 		intermediate[4095+1104:0+1104] <= intermediate[4095+1104:0+1104] + a; end
12'd1105: begin if(a[1105]==1) 
	 		intermediate[4095+1105:0+1105] <= intermediate[4095+1105:0+1105] + a; end
12'd1106: begin if(a[1106]==1) 
	 		intermediate[4095+1106:0+1106] <= intermediate[4095+1106:0+1106] + a; end
12'd1107: begin if(a[1107]==1) 
	 		intermediate[4095+1107:0+1107] <= intermediate[4095+1107:0+1107] + a; end
12'd1108: begin if(a[1108]==1) 
	 		intermediate[4095+1108:0+1108] <= intermediate[4095+1108:0+1108] + a; end
12'd1109: begin if(a[1109]==1) 
	 		intermediate[4095+1109:0+1109] <= intermediate[4095+1109:0+1109] + a; end
12'd1110: begin if(a[1110]==1) 
	 		intermediate[4095+1110:0+1110] <= intermediate[4095+1110:0+1110] + a; end
12'd1111: begin if(a[1111]==1) 
	 		intermediate[4095+1111:0+1111] <= intermediate[4095+1111:0+1111] + a; end
12'd1112: begin if(a[1112]==1) 
	 		intermediate[4095+1112:0+1112] <= intermediate[4095+1112:0+1112] + a; end
12'd1113: begin if(a[1113]==1) 
	 		intermediate[4095+1113:0+1113] <= intermediate[4095+1113:0+1113] + a; end
12'd1114: begin if(a[1114]==1) 
	 		intermediate[4095+1114:0+1114] <= intermediate[4095+1114:0+1114] + a; end
12'd1115: begin if(a[1115]==1) 
	 		intermediate[4095+1115:0+1115] <= intermediate[4095+1115:0+1115] + a; end
12'd1116: begin if(a[1116]==1) 
	 		intermediate[4095+1116:0+1116] <= intermediate[4095+1116:0+1116] + a; end
12'd1117: begin if(a[1117]==1) 
	 		intermediate[4095+1117:0+1117] <= intermediate[4095+1117:0+1117] + a; end
12'd1118: begin if(a[1118]==1) 
	 		intermediate[4095+1118:0+1118] <= intermediate[4095+1118:0+1118] + a; end
12'd1119: begin if(a[1119]==1) 
	 		intermediate[4095+1119:0+1119] <= intermediate[4095+1119:0+1119] + a; end
12'd1120: begin if(a[1120]==1) 
	 		intermediate[4095+1120:0+1120] <= intermediate[4095+1120:0+1120] + a; end
12'd1121: begin if(a[1121]==1) 
	 		intermediate[4095+1121:0+1121] <= intermediate[4095+1121:0+1121] + a; end
12'd1122: begin if(a[1122]==1) 
	 		intermediate[4095+1122:0+1122] <= intermediate[4095+1122:0+1122] + a; end
12'd1123: begin if(a[1123]==1) 
	 		intermediate[4095+1123:0+1123] <= intermediate[4095+1123:0+1123] + a; end
12'd1124: begin if(a[1124]==1) 
	 		intermediate[4095+1124:0+1124] <= intermediate[4095+1124:0+1124] + a; end
12'd1125: begin if(a[1125]==1) 
	 		intermediate[4095+1125:0+1125] <= intermediate[4095+1125:0+1125] + a; end
12'd1126: begin if(a[1126]==1) 
	 		intermediate[4095+1126:0+1126] <= intermediate[4095+1126:0+1126] + a; end
12'd1127: begin if(a[1127]==1) 
	 		intermediate[4095+1127:0+1127] <= intermediate[4095+1127:0+1127] + a; end
12'd1128: begin if(a[1128]==1) 
	 		intermediate[4095+1128:0+1128] <= intermediate[4095+1128:0+1128] + a; end
12'd1129: begin if(a[1129]==1) 
	 		intermediate[4095+1129:0+1129] <= intermediate[4095+1129:0+1129] + a; end
12'd1130: begin if(a[1130]==1) 
	 		intermediate[4095+1130:0+1130] <= intermediate[4095+1130:0+1130] + a; end
12'd1131: begin if(a[1131]==1) 
	 		intermediate[4095+1131:0+1131] <= intermediate[4095+1131:0+1131] + a; end
12'd1132: begin if(a[1132]==1) 
	 		intermediate[4095+1132:0+1132] <= intermediate[4095+1132:0+1132] + a; end
12'd1133: begin if(a[1133]==1) 
	 		intermediate[4095+1133:0+1133] <= intermediate[4095+1133:0+1133] + a; end
12'd1134: begin if(a[1134]==1) 
	 		intermediate[4095+1134:0+1134] <= intermediate[4095+1134:0+1134] + a; end
12'd1135: begin if(a[1135]==1) 
	 		intermediate[4095+1135:0+1135] <= intermediate[4095+1135:0+1135] + a; end
12'd1136: begin if(a[1136]==1) 
	 		intermediate[4095+1136:0+1136] <= intermediate[4095+1136:0+1136] + a; end
12'd1137: begin if(a[1137]==1) 
	 		intermediate[4095+1137:0+1137] <= intermediate[4095+1137:0+1137] + a; end
12'd1138: begin if(a[1138]==1) 
	 		intermediate[4095+1138:0+1138] <= intermediate[4095+1138:0+1138] + a; end
12'd1139: begin if(a[1139]==1) 
	 		intermediate[4095+1139:0+1139] <= intermediate[4095+1139:0+1139] + a; end
12'd1140: begin if(a[1140]==1) 
	 		intermediate[4095+1140:0+1140] <= intermediate[4095+1140:0+1140] + a; end
12'd1141: begin if(a[1141]==1) 
	 		intermediate[4095+1141:0+1141] <= intermediate[4095+1141:0+1141] + a; end
12'd1142: begin if(a[1142]==1) 
	 		intermediate[4095+1142:0+1142] <= intermediate[4095+1142:0+1142] + a; end
12'd1143: begin if(a[1143]==1) 
	 		intermediate[4095+1143:0+1143] <= intermediate[4095+1143:0+1143] + a; end
12'd1144: begin if(a[1144]==1) 
	 		intermediate[4095+1144:0+1144] <= intermediate[4095+1144:0+1144] + a; end
12'd1145: begin if(a[1145]==1) 
	 		intermediate[4095+1145:0+1145] <= intermediate[4095+1145:0+1145] + a; end
12'd1146: begin if(a[1146]==1) 
	 		intermediate[4095+1146:0+1146] <= intermediate[4095+1146:0+1146] + a; end
12'd1147: begin if(a[1147]==1) 
	 		intermediate[4095+1147:0+1147] <= intermediate[4095+1147:0+1147] + a; end
12'd1148: begin if(a[1148]==1) 
	 		intermediate[4095+1148:0+1148] <= intermediate[4095+1148:0+1148] + a; end
12'd1149: begin if(a[1149]==1) 
	 		intermediate[4095+1149:0+1149] <= intermediate[4095+1149:0+1149] + a; end
12'd1150: begin if(a[1150]==1) 
	 		intermediate[4095+1150:0+1150] <= intermediate[4095+1150:0+1150] + a; end
12'd1151: begin if(a[1151]==1) 
	 		intermediate[4095+1151:0+1151] <= intermediate[4095+1151:0+1151] + a; end
12'd1152: begin if(a[1152]==1) 
	 		intermediate[4095+1152:0+1152] <= intermediate[4095+1152:0+1152] + a; end
12'd1153: begin if(a[1153]==1) 
	 		intermediate[4095+1153:0+1153] <= intermediate[4095+1153:0+1153] + a; end
12'd1154: begin if(a[1154]==1) 
	 		intermediate[4095+1154:0+1154] <= intermediate[4095+1154:0+1154] + a; end
12'd1155: begin if(a[1155]==1) 
	 		intermediate[4095+1155:0+1155] <= intermediate[4095+1155:0+1155] + a; end
12'd1156: begin if(a[1156]==1) 
	 		intermediate[4095+1156:0+1156] <= intermediate[4095+1156:0+1156] + a; end
12'd1157: begin if(a[1157]==1) 
	 		intermediate[4095+1157:0+1157] <= intermediate[4095+1157:0+1157] + a; end
12'd1158: begin if(a[1158]==1) 
	 		intermediate[4095+1158:0+1158] <= intermediate[4095+1158:0+1158] + a; end
12'd1159: begin if(a[1159]==1) 
	 		intermediate[4095+1159:0+1159] <= intermediate[4095+1159:0+1159] + a; end
12'd1160: begin if(a[1160]==1) 
	 		intermediate[4095+1160:0+1160] <= intermediate[4095+1160:0+1160] + a; end
12'd1161: begin if(a[1161]==1) 
	 		intermediate[4095+1161:0+1161] <= intermediate[4095+1161:0+1161] + a; end
12'd1162: begin if(a[1162]==1) 
	 		intermediate[4095+1162:0+1162] <= intermediate[4095+1162:0+1162] + a; end
12'd1163: begin if(a[1163]==1) 
	 		intermediate[4095+1163:0+1163] <= intermediate[4095+1163:0+1163] + a; end
12'd1164: begin if(a[1164]==1) 
	 		intermediate[4095+1164:0+1164] <= intermediate[4095+1164:0+1164] + a; end
12'd1165: begin if(a[1165]==1) 
	 		intermediate[4095+1165:0+1165] <= intermediate[4095+1165:0+1165] + a; end
12'd1166: begin if(a[1166]==1) 
	 		intermediate[4095+1166:0+1166] <= intermediate[4095+1166:0+1166] + a; end
12'd1167: begin if(a[1167]==1) 
	 		intermediate[4095+1167:0+1167] <= intermediate[4095+1167:0+1167] + a; end
12'd1168: begin if(a[1168]==1) 
	 		intermediate[4095+1168:0+1168] <= intermediate[4095+1168:0+1168] + a; end
12'd1169: begin if(a[1169]==1) 
	 		intermediate[4095+1169:0+1169] <= intermediate[4095+1169:0+1169] + a; end
12'd1170: begin if(a[1170]==1) 
	 		intermediate[4095+1170:0+1170] <= intermediate[4095+1170:0+1170] + a; end
12'd1171: begin if(a[1171]==1) 
	 		intermediate[4095+1171:0+1171] <= intermediate[4095+1171:0+1171] + a; end
12'd1172: begin if(a[1172]==1) 
	 		intermediate[4095+1172:0+1172] <= intermediate[4095+1172:0+1172] + a; end
12'd1173: begin if(a[1173]==1) 
	 		intermediate[4095+1173:0+1173] <= intermediate[4095+1173:0+1173] + a; end
12'd1174: begin if(a[1174]==1) 
	 		intermediate[4095+1174:0+1174] <= intermediate[4095+1174:0+1174] + a; end
12'd1175: begin if(a[1175]==1) 
	 		intermediate[4095+1175:0+1175] <= intermediate[4095+1175:0+1175] + a; end
12'd1176: begin if(a[1176]==1) 
	 		intermediate[4095+1176:0+1176] <= intermediate[4095+1176:0+1176] + a; end
12'd1177: begin if(a[1177]==1) 
	 		intermediate[4095+1177:0+1177] <= intermediate[4095+1177:0+1177] + a; end
12'd1178: begin if(a[1178]==1) 
	 		intermediate[4095+1178:0+1178] <= intermediate[4095+1178:0+1178] + a; end
12'd1179: begin if(a[1179]==1) 
	 		intermediate[4095+1179:0+1179] <= intermediate[4095+1179:0+1179] + a; end
12'd1180: begin if(a[1180]==1) 
	 		intermediate[4095+1180:0+1180] <= intermediate[4095+1180:0+1180] + a; end
12'd1181: begin if(a[1181]==1) 
	 		intermediate[4095+1181:0+1181] <= intermediate[4095+1181:0+1181] + a; end
12'd1182: begin if(a[1182]==1) 
	 		intermediate[4095+1182:0+1182] <= intermediate[4095+1182:0+1182] + a; end
12'd1183: begin if(a[1183]==1) 
	 		intermediate[4095+1183:0+1183] <= intermediate[4095+1183:0+1183] + a; end
12'd1184: begin if(a[1184]==1) 
	 		intermediate[4095+1184:0+1184] <= intermediate[4095+1184:0+1184] + a; end
12'd1185: begin if(a[1185]==1) 
	 		intermediate[4095+1185:0+1185] <= intermediate[4095+1185:0+1185] + a; end
12'd1186: begin if(a[1186]==1) 
	 		intermediate[4095+1186:0+1186] <= intermediate[4095+1186:0+1186] + a; end
12'd1187: begin if(a[1187]==1) 
	 		intermediate[4095+1187:0+1187] <= intermediate[4095+1187:0+1187] + a; end
12'd1188: begin if(a[1188]==1) 
	 		intermediate[4095+1188:0+1188] <= intermediate[4095+1188:0+1188] + a; end
12'd1189: begin if(a[1189]==1) 
	 		intermediate[4095+1189:0+1189] <= intermediate[4095+1189:0+1189] + a; end
12'd1190: begin if(a[1190]==1) 
	 		intermediate[4095+1190:0+1190] <= intermediate[4095+1190:0+1190] + a; end
12'd1191: begin if(a[1191]==1) 
	 		intermediate[4095+1191:0+1191] <= intermediate[4095+1191:0+1191] + a; end
12'd1192: begin if(a[1192]==1) 
	 		intermediate[4095+1192:0+1192] <= intermediate[4095+1192:0+1192] + a; end
12'd1193: begin if(a[1193]==1) 
	 		intermediate[4095+1193:0+1193] <= intermediate[4095+1193:0+1193] + a; end
12'd1194: begin if(a[1194]==1) 
	 		intermediate[4095+1194:0+1194] <= intermediate[4095+1194:0+1194] + a; end
12'd1195: begin if(a[1195]==1) 
	 		intermediate[4095+1195:0+1195] <= intermediate[4095+1195:0+1195] + a; end
12'd1196: begin if(a[1196]==1) 
	 		intermediate[4095+1196:0+1196] <= intermediate[4095+1196:0+1196] + a; end
12'd1197: begin if(a[1197]==1) 
	 		intermediate[4095+1197:0+1197] <= intermediate[4095+1197:0+1197] + a; end
12'd1198: begin if(a[1198]==1) 
	 		intermediate[4095+1198:0+1198] <= intermediate[4095+1198:0+1198] + a; end
12'd1199: begin if(a[1199]==1) 
	 		intermediate[4095+1199:0+1199] <= intermediate[4095+1199:0+1199] + a; end
12'd1200: begin if(a[1200]==1) 
	 		intermediate[4095+1200:0+1200] <= intermediate[4095+1200:0+1200] + a; end
12'd1201: begin if(a[1201]==1) 
	 		intermediate[4095+1201:0+1201] <= intermediate[4095+1201:0+1201] + a; end
12'd1202: begin if(a[1202]==1) 
	 		intermediate[4095+1202:0+1202] <= intermediate[4095+1202:0+1202] + a; end
12'd1203: begin if(a[1203]==1) 
	 		intermediate[4095+1203:0+1203] <= intermediate[4095+1203:0+1203] + a; end
12'd1204: begin if(a[1204]==1) 
	 		intermediate[4095+1204:0+1204] <= intermediate[4095+1204:0+1204] + a; end
12'd1205: begin if(a[1205]==1) 
	 		intermediate[4095+1205:0+1205] <= intermediate[4095+1205:0+1205] + a; end
12'd1206: begin if(a[1206]==1) 
	 		intermediate[4095+1206:0+1206] <= intermediate[4095+1206:0+1206] + a; end
12'd1207: begin if(a[1207]==1) 
	 		intermediate[4095+1207:0+1207] <= intermediate[4095+1207:0+1207] + a; end
12'd1208: begin if(a[1208]==1) 
	 		intermediate[4095+1208:0+1208] <= intermediate[4095+1208:0+1208] + a; end
12'd1209: begin if(a[1209]==1) 
	 		intermediate[4095+1209:0+1209] <= intermediate[4095+1209:0+1209] + a; end
12'd1210: begin if(a[1210]==1) 
	 		intermediate[4095+1210:0+1210] <= intermediate[4095+1210:0+1210] + a; end
12'd1211: begin if(a[1211]==1) 
	 		intermediate[4095+1211:0+1211] <= intermediate[4095+1211:0+1211] + a; end
12'd1212: begin if(a[1212]==1) 
	 		intermediate[4095+1212:0+1212] <= intermediate[4095+1212:0+1212] + a; end
12'd1213: begin if(a[1213]==1) 
	 		intermediate[4095+1213:0+1213] <= intermediate[4095+1213:0+1213] + a; end
12'd1214: begin if(a[1214]==1) 
	 		intermediate[4095+1214:0+1214] <= intermediate[4095+1214:0+1214] + a; end
12'd1215: begin if(a[1215]==1) 
	 		intermediate[4095+1215:0+1215] <= intermediate[4095+1215:0+1215] + a; end
12'd1216: begin if(a[1216]==1) 
	 		intermediate[4095+1216:0+1216] <= intermediate[4095+1216:0+1216] + a; end
12'd1217: begin if(a[1217]==1) 
	 		intermediate[4095+1217:0+1217] <= intermediate[4095+1217:0+1217] + a; end
12'd1218: begin if(a[1218]==1) 
	 		intermediate[4095+1218:0+1218] <= intermediate[4095+1218:0+1218] + a; end
12'd1219: begin if(a[1219]==1) 
	 		intermediate[4095+1219:0+1219] <= intermediate[4095+1219:0+1219] + a; end
12'd1220: begin if(a[1220]==1) 
	 		intermediate[4095+1220:0+1220] <= intermediate[4095+1220:0+1220] + a; end
12'd1221: begin if(a[1221]==1) 
	 		intermediate[4095+1221:0+1221] <= intermediate[4095+1221:0+1221] + a; end
12'd1222: begin if(a[1222]==1) 
	 		intermediate[4095+1222:0+1222] <= intermediate[4095+1222:0+1222] + a; end
12'd1223: begin if(a[1223]==1) 
	 		intermediate[4095+1223:0+1223] <= intermediate[4095+1223:0+1223] + a; end
12'd1224: begin if(a[1224]==1) 
	 		intermediate[4095+1224:0+1224] <= intermediate[4095+1224:0+1224] + a; end
12'd1225: begin if(a[1225]==1) 
	 		intermediate[4095+1225:0+1225] <= intermediate[4095+1225:0+1225] + a; end
12'd1226: begin if(a[1226]==1) 
	 		intermediate[4095+1226:0+1226] <= intermediate[4095+1226:0+1226] + a; end
12'd1227: begin if(a[1227]==1) 
	 		intermediate[4095+1227:0+1227] <= intermediate[4095+1227:0+1227] + a; end
12'd1228: begin if(a[1228]==1) 
	 		intermediate[4095+1228:0+1228] <= intermediate[4095+1228:0+1228] + a; end
12'd1229: begin if(a[1229]==1) 
	 		intermediate[4095+1229:0+1229] <= intermediate[4095+1229:0+1229] + a; end
12'd1230: begin if(a[1230]==1) 
	 		intermediate[4095+1230:0+1230] <= intermediate[4095+1230:0+1230] + a; end
12'd1231: begin if(a[1231]==1) 
	 		intermediate[4095+1231:0+1231] <= intermediate[4095+1231:0+1231] + a; end
12'd1232: begin if(a[1232]==1) 
	 		intermediate[4095+1232:0+1232] <= intermediate[4095+1232:0+1232] + a; end
12'd1233: begin if(a[1233]==1) 
	 		intermediate[4095+1233:0+1233] <= intermediate[4095+1233:0+1233] + a; end
12'd1234: begin if(a[1234]==1) 
	 		intermediate[4095+1234:0+1234] <= intermediate[4095+1234:0+1234] + a; end
12'd1235: begin if(a[1235]==1) 
	 		intermediate[4095+1235:0+1235] <= intermediate[4095+1235:0+1235] + a; end
12'd1236: begin if(a[1236]==1) 
	 		intermediate[4095+1236:0+1236] <= intermediate[4095+1236:0+1236] + a; end
12'd1237: begin if(a[1237]==1) 
	 		intermediate[4095+1237:0+1237] <= intermediate[4095+1237:0+1237] + a; end
12'd1238: begin if(a[1238]==1) 
	 		intermediate[4095+1238:0+1238] <= intermediate[4095+1238:0+1238] + a; end
12'd1239: begin if(a[1239]==1) 
	 		intermediate[4095+1239:0+1239] <= intermediate[4095+1239:0+1239] + a; end
12'd1240: begin if(a[1240]==1) 
	 		intermediate[4095+1240:0+1240] <= intermediate[4095+1240:0+1240] + a; end
12'd1241: begin if(a[1241]==1) 
	 		intermediate[4095+1241:0+1241] <= intermediate[4095+1241:0+1241] + a; end
12'd1242: begin if(a[1242]==1) 
	 		intermediate[4095+1242:0+1242] <= intermediate[4095+1242:0+1242] + a; end
12'd1243: begin if(a[1243]==1) 
	 		intermediate[4095+1243:0+1243] <= intermediate[4095+1243:0+1243] + a; end
12'd1244: begin if(a[1244]==1) 
	 		intermediate[4095+1244:0+1244] <= intermediate[4095+1244:0+1244] + a; end
12'd1245: begin if(a[1245]==1) 
	 		intermediate[4095+1245:0+1245] <= intermediate[4095+1245:0+1245] + a; end
12'd1246: begin if(a[1246]==1) 
	 		intermediate[4095+1246:0+1246] <= intermediate[4095+1246:0+1246] + a; end
12'd1247: begin if(a[1247]==1) 
	 		intermediate[4095+1247:0+1247] <= intermediate[4095+1247:0+1247] + a; end
12'd1248: begin if(a[1248]==1) 
	 		intermediate[4095+1248:0+1248] <= intermediate[4095+1248:0+1248] + a; end
12'd1249: begin if(a[1249]==1) 
	 		intermediate[4095+1249:0+1249] <= intermediate[4095+1249:0+1249] + a; end
12'd1250: begin if(a[1250]==1) 
	 		intermediate[4095+1250:0+1250] <= intermediate[4095+1250:0+1250] + a; end
12'd1251: begin if(a[1251]==1) 
	 		intermediate[4095+1251:0+1251] <= intermediate[4095+1251:0+1251] + a; end
12'd1252: begin if(a[1252]==1) 
	 		intermediate[4095+1252:0+1252] <= intermediate[4095+1252:0+1252] + a; end
12'd1253: begin if(a[1253]==1) 
	 		intermediate[4095+1253:0+1253] <= intermediate[4095+1253:0+1253] + a; end
12'd1254: begin if(a[1254]==1) 
	 		intermediate[4095+1254:0+1254] <= intermediate[4095+1254:0+1254] + a; end
12'd1255: begin if(a[1255]==1) 
	 		intermediate[4095+1255:0+1255] <= intermediate[4095+1255:0+1255] + a; end
12'd1256: begin if(a[1256]==1) 
	 		intermediate[4095+1256:0+1256] <= intermediate[4095+1256:0+1256] + a; end
12'd1257: begin if(a[1257]==1) 
	 		intermediate[4095+1257:0+1257] <= intermediate[4095+1257:0+1257] + a; end
12'd1258: begin if(a[1258]==1) 
	 		intermediate[4095+1258:0+1258] <= intermediate[4095+1258:0+1258] + a; end
12'd1259: begin if(a[1259]==1) 
	 		intermediate[4095+1259:0+1259] <= intermediate[4095+1259:0+1259] + a; end
12'd1260: begin if(a[1260]==1) 
	 		intermediate[4095+1260:0+1260] <= intermediate[4095+1260:0+1260] + a; end
12'd1261: begin if(a[1261]==1) 
	 		intermediate[4095+1261:0+1261] <= intermediate[4095+1261:0+1261] + a; end
12'd1262: begin if(a[1262]==1) 
	 		intermediate[4095+1262:0+1262] <= intermediate[4095+1262:0+1262] + a; end
12'd1263: begin if(a[1263]==1) 
	 		intermediate[4095+1263:0+1263] <= intermediate[4095+1263:0+1263] + a; end
12'd1264: begin if(a[1264]==1) 
	 		intermediate[4095+1264:0+1264] <= intermediate[4095+1264:0+1264] + a; end
12'd1265: begin if(a[1265]==1) 
	 		intermediate[4095+1265:0+1265] <= intermediate[4095+1265:0+1265] + a; end
12'd1266: begin if(a[1266]==1) 
	 		intermediate[4095+1266:0+1266] <= intermediate[4095+1266:0+1266] + a; end
12'd1267: begin if(a[1267]==1) 
	 		intermediate[4095+1267:0+1267] <= intermediate[4095+1267:0+1267] + a; end
12'd1268: begin if(a[1268]==1) 
	 		intermediate[4095+1268:0+1268] <= intermediate[4095+1268:0+1268] + a; end
12'd1269: begin if(a[1269]==1) 
	 		intermediate[4095+1269:0+1269] <= intermediate[4095+1269:0+1269] + a; end
12'd1270: begin if(a[1270]==1) 
	 		intermediate[4095+1270:0+1270] <= intermediate[4095+1270:0+1270] + a; end
12'd1271: begin if(a[1271]==1) 
	 		intermediate[4095+1271:0+1271] <= intermediate[4095+1271:0+1271] + a; end
12'd1272: begin if(a[1272]==1) 
	 		intermediate[4095+1272:0+1272] <= intermediate[4095+1272:0+1272] + a; end
12'd1273: begin if(a[1273]==1) 
	 		intermediate[4095+1273:0+1273] <= intermediate[4095+1273:0+1273] + a; end
12'd1274: begin if(a[1274]==1) 
	 		intermediate[4095+1274:0+1274] <= intermediate[4095+1274:0+1274] + a; end
12'd1275: begin if(a[1275]==1) 
	 		intermediate[4095+1275:0+1275] <= intermediate[4095+1275:0+1275] + a; end
12'd1276: begin if(a[1276]==1) 
	 		intermediate[4095+1276:0+1276] <= intermediate[4095+1276:0+1276] + a; end
12'd1277: begin if(a[1277]==1) 
	 		intermediate[4095+1277:0+1277] <= intermediate[4095+1277:0+1277] + a; end
12'd1278: begin if(a[1278]==1) 
	 		intermediate[4095+1278:0+1278] <= intermediate[4095+1278:0+1278] + a; end
12'd1279: begin if(a[1279]==1) 
	 		intermediate[4095+1279:0+1279] <= intermediate[4095+1279:0+1279] + a; end
12'd1280: begin if(a[1280]==1) 
	 		intermediate[4095+1280:0+1280] <= intermediate[4095+1280:0+1280] + a; end
12'd1281: begin if(a[1281]==1) 
	 		intermediate[4095+1281:0+1281] <= intermediate[4095+1281:0+1281] + a; end
12'd1282: begin if(a[1282]==1) 
	 		intermediate[4095+1282:0+1282] <= intermediate[4095+1282:0+1282] + a; end
12'd1283: begin if(a[1283]==1) 
	 		intermediate[4095+1283:0+1283] <= intermediate[4095+1283:0+1283] + a; end
12'd1284: begin if(a[1284]==1) 
	 		intermediate[4095+1284:0+1284] <= intermediate[4095+1284:0+1284] + a; end
12'd1285: begin if(a[1285]==1) 
	 		intermediate[4095+1285:0+1285] <= intermediate[4095+1285:0+1285] + a; end
12'd1286: begin if(a[1286]==1) 
	 		intermediate[4095+1286:0+1286] <= intermediate[4095+1286:0+1286] + a; end
12'd1287: begin if(a[1287]==1) 
	 		intermediate[4095+1287:0+1287] <= intermediate[4095+1287:0+1287] + a; end
12'd1288: begin if(a[1288]==1) 
	 		intermediate[4095+1288:0+1288] <= intermediate[4095+1288:0+1288] + a; end
12'd1289: begin if(a[1289]==1) 
	 		intermediate[4095+1289:0+1289] <= intermediate[4095+1289:0+1289] + a; end
12'd1290: begin if(a[1290]==1) 
	 		intermediate[4095+1290:0+1290] <= intermediate[4095+1290:0+1290] + a; end
12'd1291: begin if(a[1291]==1) 
	 		intermediate[4095+1291:0+1291] <= intermediate[4095+1291:0+1291] + a; end
12'd1292: begin if(a[1292]==1) 
	 		intermediate[4095+1292:0+1292] <= intermediate[4095+1292:0+1292] + a; end
12'd1293: begin if(a[1293]==1) 
	 		intermediate[4095+1293:0+1293] <= intermediate[4095+1293:0+1293] + a; end
12'd1294: begin if(a[1294]==1) 
	 		intermediate[4095+1294:0+1294] <= intermediate[4095+1294:0+1294] + a; end
12'd1295: begin if(a[1295]==1) 
	 		intermediate[4095+1295:0+1295] <= intermediate[4095+1295:0+1295] + a; end
12'd1296: begin if(a[1296]==1) 
	 		intermediate[4095+1296:0+1296] <= intermediate[4095+1296:0+1296] + a; end
12'd1297: begin if(a[1297]==1) 
	 		intermediate[4095+1297:0+1297] <= intermediate[4095+1297:0+1297] + a; end
12'd1298: begin if(a[1298]==1) 
	 		intermediate[4095+1298:0+1298] <= intermediate[4095+1298:0+1298] + a; end
12'd1299: begin if(a[1299]==1) 
	 		intermediate[4095+1299:0+1299] <= intermediate[4095+1299:0+1299] + a; end
12'd1300: begin if(a[1300]==1) 
	 		intermediate[4095+1300:0+1300] <= intermediate[4095+1300:0+1300] + a; end
12'd1301: begin if(a[1301]==1) 
	 		intermediate[4095+1301:0+1301] <= intermediate[4095+1301:0+1301] + a; end
12'd1302: begin if(a[1302]==1) 
	 		intermediate[4095+1302:0+1302] <= intermediate[4095+1302:0+1302] + a; end
12'd1303: begin if(a[1303]==1) 
	 		intermediate[4095+1303:0+1303] <= intermediate[4095+1303:0+1303] + a; end
12'd1304: begin if(a[1304]==1) 
	 		intermediate[4095+1304:0+1304] <= intermediate[4095+1304:0+1304] + a; end
12'd1305: begin if(a[1305]==1) 
	 		intermediate[4095+1305:0+1305] <= intermediate[4095+1305:0+1305] + a; end
12'd1306: begin if(a[1306]==1) 
	 		intermediate[4095+1306:0+1306] <= intermediate[4095+1306:0+1306] + a; end
12'd1307: begin if(a[1307]==1) 
	 		intermediate[4095+1307:0+1307] <= intermediate[4095+1307:0+1307] + a; end
12'd1308: begin if(a[1308]==1) 
	 		intermediate[4095+1308:0+1308] <= intermediate[4095+1308:0+1308] + a; end
12'd1309: begin if(a[1309]==1) 
	 		intermediate[4095+1309:0+1309] <= intermediate[4095+1309:0+1309] + a; end
12'd1310: begin if(a[1310]==1) 
	 		intermediate[4095+1310:0+1310] <= intermediate[4095+1310:0+1310] + a; end
12'd1311: begin if(a[1311]==1) 
	 		intermediate[4095+1311:0+1311] <= intermediate[4095+1311:0+1311] + a; end
12'd1312: begin if(a[1312]==1) 
	 		intermediate[4095+1312:0+1312] <= intermediate[4095+1312:0+1312] + a; end
12'd1313: begin if(a[1313]==1) 
	 		intermediate[4095+1313:0+1313] <= intermediate[4095+1313:0+1313] + a; end
12'd1314: begin if(a[1314]==1) 
	 		intermediate[4095+1314:0+1314] <= intermediate[4095+1314:0+1314] + a; end
12'd1315: begin if(a[1315]==1) 
	 		intermediate[4095+1315:0+1315] <= intermediate[4095+1315:0+1315] + a; end
12'd1316: begin if(a[1316]==1) 
	 		intermediate[4095+1316:0+1316] <= intermediate[4095+1316:0+1316] + a; end
12'd1317: begin if(a[1317]==1) 
	 		intermediate[4095+1317:0+1317] <= intermediate[4095+1317:0+1317] + a; end
12'd1318: begin if(a[1318]==1) 
	 		intermediate[4095+1318:0+1318] <= intermediate[4095+1318:0+1318] + a; end
12'd1319: begin if(a[1319]==1) 
	 		intermediate[4095+1319:0+1319] <= intermediate[4095+1319:0+1319] + a; end
12'd1320: begin if(a[1320]==1) 
	 		intermediate[4095+1320:0+1320] <= intermediate[4095+1320:0+1320] + a; end
12'd1321: begin if(a[1321]==1) 
	 		intermediate[4095+1321:0+1321] <= intermediate[4095+1321:0+1321] + a; end
12'd1322: begin if(a[1322]==1) 
	 		intermediate[4095+1322:0+1322] <= intermediate[4095+1322:0+1322] + a; end
12'd1323: begin if(a[1323]==1) 
	 		intermediate[4095+1323:0+1323] <= intermediate[4095+1323:0+1323] + a; end
12'd1324: begin if(a[1324]==1) 
	 		intermediate[4095+1324:0+1324] <= intermediate[4095+1324:0+1324] + a; end
12'd1325: begin if(a[1325]==1) 
	 		intermediate[4095+1325:0+1325] <= intermediate[4095+1325:0+1325] + a; end
12'd1326: begin if(a[1326]==1) 
	 		intermediate[4095+1326:0+1326] <= intermediate[4095+1326:0+1326] + a; end
12'd1327: begin if(a[1327]==1) 
	 		intermediate[4095+1327:0+1327] <= intermediate[4095+1327:0+1327] + a; end
12'd1328: begin if(a[1328]==1) 
	 		intermediate[4095+1328:0+1328] <= intermediate[4095+1328:0+1328] + a; end
12'd1329: begin if(a[1329]==1) 
	 		intermediate[4095+1329:0+1329] <= intermediate[4095+1329:0+1329] + a; end
12'd1330: begin if(a[1330]==1) 
	 		intermediate[4095+1330:0+1330] <= intermediate[4095+1330:0+1330] + a; end
12'd1331: begin if(a[1331]==1) 
	 		intermediate[4095+1331:0+1331] <= intermediate[4095+1331:0+1331] + a; end
12'd1332: begin if(a[1332]==1) 
	 		intermediate[4095+1332:0+1332] <= intermediate[4095+1332:0+1332] + a; end
12'd1333: begin if(a[1333]==1) 
	 		intermediate[4095+1333:0+1333] <= intermediate[4095+1333:0+1333] + a; end
12'd1334: begin if(a[1334]==1) 
	 		intermediate[4095+1334:0+1334] <= intermediate[4095+1334:0+1334] + a; end
12'd1335: begin if(a[1335]==1) 
	 		intermediate[4095+1335:0+1335] <= intermediate[4095+1335:0+1335] + a; end
12'd1336: begin if(a[1336]==1) 
	 		intermediate[4095+1336:0+1336] <= intermediate[4095+1336:0+1336] + a; end
12'd1337: begin if(a[1337]==1) 
	 		intermediate[4095+1337:0+1337] <= intermediate[4095+1337:0+1337] + a; end
12'd1338: begin if(a[1338]==1) 
	 		intermediate[4095+1338:0+1338] <= intermediate[4095+1338:0+1338] + a; end
12'd1339: begin if(a[1339]==1) 
	 		intermediate[4095+1339:0+1339] <= intermediate[4095+1339:0+1339] + a; end
12'd1340: begin if(a[1340]==1) 
	 		intermediate[4095+1340:0+1340] <= intermediate[4095+1340:0+1340] + a; end
12'd1341: begin if(a[1341]==1) 
	 		intermediate[4095+1341:0+1341] <= intermediate[4095+1341:0+1341] + a; end
12'd1342: begin if(a[1342]==1) 
	 		intermediate[4095+1342:0+1342] <= intermediate[4095+1342:0+1342] + a; end
12'd1343: begin if(a[1343]==1) 
	 		intermediate[4095+1343:0+1343] <= intermediate[4095+1343:0+1343] + a; end
12'd1344: begin if(a[1344]==1) 
	 		intermediate[4095+1344:0+1344] <= intermediate[4095+1344:0+1344] + a; end
12'd1345: begin if(a[1345]==1) 
	 		intermediate[4095+1345:0+1345] <= intermediate[4095+1345:0+1345] + a; end
12'd1346: begin if(a[1346]==1) 
	 		intermediate[4095+1346:0+1346] <= intermediate[4095+1346:0+1346] + a; end
12'd1347: begin if(a[1347]==1) 
	 		intermediate[4095+1347:0+1347] <= intermediate[4095+1347:0+1347] + a; end
12'd1348: begin if(a[1348]==1) 
	 		intermediate[4095+1348:0+1348] <= intermediate[4095+1348:0+1348] + a; end
12'd1349: begin if(a[1349]==1) 
	 		intermediate[4095+1349:0+1349] <= intermediate[4095+1349:0+1349] + a; end
12'd1350: begin if(a[1350]==1) 
	 		intermediate[4095+1350:0+1350] <= intermediate[4095+1350:0+1350] + a; end
12'd1351: begin if(a[1351]==1) 
	 		intermediate[4095+1351:0+1351] <= intermediate[4095+1351:0+1351] + a; end
12'd1352: begin if(a[1352]==1) 
	 		intermediate[4095+1352:0+1352] <= intermediate[4095+1352:0+1352] + a; end
12'd1353: begin if(a[1353]==1) 
	 		intermediate[4095+1353:0+1353] <= intermediate[4095+1353:0+1353] + a; end
12'd1354: begin if(a[1354]==1) 
	 		intermediate[4095+1354:0+1354] <= intermediate[4095+1354:0+1354] + a; end
12'd1355: begin if(a[1355]==1) 
	 		intermediate[4095+1355:0+1355] <= intermediate[4095+1355:0+1355] + a; end
12'd1356: begin if(a[1356]==1) 
	 		intermediate[4095+1356:0+1356] <= intermediate[4095+1356:0+1356] + a; end
12'd1357: begin if(a[1357]==1) 
	 		intermediate[4095+1357:0+1357] <= intermediate[4095+1357:0+1357] + a; end
12'd1358: begin if(a[1358]==1) 
	 		intermediate[4095+1358:0+1358] <= intermediate[4095+1358:0+1358] + a; end
12'd1359: begin if(a[1359]==1) 
	 		intermediate[4095+1359:0+1359] <= intermediate[4095+1359:0+1359] + a; end
12'd1360: begin if(a[1360]==1) 
	 		intermediate[4095+1360:0+1360] <= intermediate[4095+1360:0+1360] + a; end
12'd1361: begin if(a[1361]==1) 
	 		intermediate[4095+1361:0+1361] <= intermediate[4095+1361:0+1361] + a; end
12'd1362: begin if(a[1362]==1) 
	 		intermediate[4095+1362:0+1362] <= intermediate[4095+1362:0+1362] + a; end
12'd1363: begin if(a[1363]==1) 
	 		intermediate[4095+1363:0+1363] <= intermediate[4095+1363:0+1363] + a; end
12'd1364: begin if(a[1364]==1) 
	 		intermediate[4095+1364:0+1364] <= intermediate[4095+1364:0+1364] + a; end
12'd1365: begin if(a[1365]==1) 
	 		intermediate[4095+1365:0+1365] <= intermediate[4095+1365:0+1365] + a; end
12'd1366: begin if(a[1366]==1) 
	 		intermediate[4095+1366:0+1366] <= intermediate[4095+1366:0+1366] + a; end
12'd1367: begin if(a[1367]==1) 
	 		intermediate[4095+1367:0+1367] <= intermediate[4095+1367:0+1367] + a; end
12'd1368: begin if(a[1368]==1) 
	 		intermediate[4095+1368:0+1368] <= intermediate[4095+1368:0+1368] + a; end
12'd1369: begin if(a[1369]==1) 
	 		intermediate[4095+1369:0+1369] <= intermediate[4095+1369:0+1369] + a; end
12'd1370: begin if(a[1370]==1) 
	 		intermediate[4095+1370:0+1370] <= intermediate[4095+1370:0+1370] + a; end
12'd1371: begin if(a[1371]==1) 
	 		intermediate[4095+1371:0+1371] <= intermediate[4095+1371:0+1371] + a; end
12'd1372: begin if(a[1372]==1) 
	 		intermediate[4095+1372:0+1372] <= intermediate[4095+1372:0+1372] + a; end
12'd1373: begin if(a[1373]==1) 
	 		intermediate[4095+1373:0+1373] <= intermediate[4095+1373:0+1373] + a; end
12'd1374: begin if(a[1374]==1) 
	 		intermediate[4095+1374:0+1374] <= intermediate[4095+1374:0+1374] + a; end
12'd1375: begin if(a[1375]==1) 
	 		intermediate[4095+1375:0+1375] <= intermediate[4095+1375:0+1375] + a; end
12'd1376: begin if(a[1376]==1) 
	 		intermediate[4095+1376:0+1376] <= intermediate[4095+1376:0+1376] + a; end
12'd1377: begin if(a[1377]==1) 
	 		intermediate[4095+1377:0+1377] <= intermediate[4095+1377:0+1377] + a; end
12'd1378: begin if(a[1378]==1) 
	 		intermediate[4095+1378:0+1378] <= intermediate[4095+1378:0+1378] + a; end
12'd1379: begin if(a[1379]==1) 
	 		intermediate[4095+1379:0+1379] <= intermediate[4095+1379:0+1379] + a; end
12'd1380: begin if(a[1380]==1) 
	 		intermediate[4095+1380:0+1380] <= intermediate[4095+1380:0+1380] + a; end
12'd1381: begin if(a[1381]==1) 
	 		intermediate[4095+1381:0+1381] <= intermediate[4095+1381:0+1381] + a; end
12'd1382: begin if(a[1382]==1) 
	 		intermediate[4095+1382:0+1382] <= intermediate[4095+1382:0+1382] + a; end
12'd1383: begin if(a[1383]==1) 
	 		intermediate[4095+1383:0+1383] <= intermediate[4095+1383:0+1383] + a; end
12'd1384: begin if(a[1384]==1) 
	 		intermediate[4095+1384:0+1384] <= intermediate[4095+1384:0+1384] + a; end
12'd1385: begin if(a[1385]==1) 
	 		intermediate[4095+1385:0+1385] <= intermediate[4095+1385:0+1385] + a; end
12'd1386: begin if(a[1386]==1) 
	 		intermediate[4095+1386:0+1386] <= intermediate[4095+1386:0+1386] + a; end
12'd1387: begin if(a[1387]==1) 
	 		intermediate[4095+1387:0+1387] <= intermediate[4095+1387:0+1387] + a; end
12'd1388: begin if(a[1388]==1) 
	 		intermediate[4095+1388:0+1388] <= intermediate[4095+1388:0+1388] + a; end
12'd1389: begin if(a[1389]==1) 
	 		intermediate[4095+1389:0+1389] <= intermediate[4095+1389:0+1389] + a; end
12'd1390: begin if(a[1390]==1) 
	 		intermediate[4095+1390:0+1390] <= intermediate[4095+1390:0+1390] + a; end
12'd1391: begin if(a[1391]==1) 
	 		intermediate[4095+1391:0+1391] <= intermediate[4095+1391:0+1391] + a; end
12'd1392: begin if(a[1392]==1) 
	 		intermediate[4095+1392:0+1392] <= intermediate[4095+1392:0+1392] + a; end
12'd1393: begin if(a[1393]==1) 
	 		intermediate[4095+1393:0+1393] <= intermediate[4095+1393:0+1393] + a; end
12'd1394: begin if(a[1394]==1) 
	 		intermediate[4095+1394:0+1394] <= intermediate[4095+1394:0+1394] + a; end
12'd1395: begin if(a[1395]==1) 
	 		intermediate[4095+1395:0+1395] <= intermediate[4095+1395:0+1395] + a; end
12'd1396: begin if(a[1396]==1) 
	 		intermediate[4095+1396:0+1396] <= intermediate[4095+1396:0+1396] + a; end
12'd1397: begin if(a[1397]==1) 
	 		intermediate[4095+1397:0+1397] <= intermediate[4095+1397:0+1397] + a; end
12'd1398: begin if(a[1398]==1) 
	 		intermediate[4095+1398:0+1398] <= intermediate[4095+1398:0+1398] + a; end
12'd1399: begin if(a[1399]==1) 
	 		intermediate[4095+1399:0+1399] <= intermediate[4095+1399:0+1399] + a; end
12'd1400: begin if(a[1400]==1) 
	 		intermediate[4095+1400:0+1400] <= intermediate[4095+1400:0+1400] + a; end
12'd1401: begin if(a[1401]==1) 
	 		intermediate[4095+1401:0+1401] <= intermediate[4095+1401:0+1401] + a; end
12'd1402: begin if(a[1402]==1) 
	 		intermediate[4095+1402:0+1402] <= intermediate[4095+1402:0+1402] + a; end
12'd1403: begin if(a[1403]==1) 
	 		intermediate[4095+1403:0+1403] <= intermediate[4095+1403:0+1403] + a; end
12'd1404: begin if(a[1404]==1) 
	 		intermediate[4095+1404:0+1404] <= intermediate[4095+1404:0+1404] + a; end
12'd1405: begin if(a[1405]==1) 
	 		intermediate[4095+1405:0+1405] <= intermediate[4095+1405:0+1405] + a; end
12'd1406: begin if(a[1406]==1) 
	 		intermediate[4095+1406:0+1406] <= intermediate[4095+1406:0+1406] + a; end
12'd1407: begin if(a[1407]==1) 
	 		intermediate[4095+1407:0+1407] <= intermediate[4095+1407:0+1407] + a; end
12'd1408: begin if(a[1408]==1) 
	 		intermediate[4095+1408:0+1408] <= intermediate[4095+1408:0+1408] + a; end
12'd1409: begin if(a[1409]==1) 
	 		intermediate[4095+1409:0+1409] <= intermediate[4095+1409:0+1409] + a; end
12'd1410: begin if(a[1410]==1) 
	 		intermediate[4095+1410:0+1410] <= intermediate[4095+1410:0+1410] + a; end
12'd1411: begin if(a[1411]==1) 
	 		intermediate[4095+1411:0+1411] <= intermediate[4095+1411:0+1411] + a; end
12'd1412: begin if(a[1412]==1) 
	 		intermediate[4095+1412:0+1412] <= intermediate[4095+1412:0+1412] + a; end
12'd1413: begin if(a[1413]==1) 
	 		intermediate[4095+1413:0+1413] <= intermediate[4095+1413:0+1413] + a; end
12'd1414: begin if(a[1414]==1) 
	 		intermediate[4095+1414:0+1414] <= intermediate[4095+1414:0+1414] + a; end
12'd1415: begin if(a[1415]==1) 
	 		intermediate[4095+1415:0+1415] <= intermediate[4095+1415:0+1415] + a; end
12'd1416: begin if(a[1416]==1) 
	 		intermediate[4095+1416:0+1416] <= intermediate[4095+1416:0+1416] + a; end
12'd1417: begin if(a[1417]==1) 
	 		intermediate[4095+1417:0+1417] <= intermediate[4095+1417:0+1417] + a; end
12'd1418: begin if(a[1418]==1) 
	 		intermediate[4095+1418:0+1418] <= intermediate[4095+1418:0+1418] + a; end
12'd1419: begin if(a[1419]==1) 
	 		intermediate[4095+1419:0+1419] <= intermediate[4095+1419:0+1419] + a; end
12'd1420: begin if(a[1420]==1) 
	 		intermediate[4095+1420:0+1420] <= intermediate[4095+1420:0+1420] + a; end
12'd1421: begin if(a[1421]==1) 
	 		intermediate[4095+1421:0+1421] <= intermediate[4095+1421:0+1421] + a; end
12'd1422: begin if(a[1422]==1) 
	 		intermediate[4095+1422:0+1422] <= intermediate[4095+1422:0+1422] + a; end
12'd1423: begin if(a[1423]==1) 
	 		intermediate[4095+1423:0+1423] <= intermediate[4095+1423:0+1423] + a; end
12'd1424: begin if(a[1424]==1) 
	 		intermediate[4095+1424:0+1424] <= intermediate[4095+1424:0+1424] + a; end
12'd1425: begin if(a[1425]==1) 
	 		intermediate[4095+1425:0+1425] <= intermediate[4095+1425:0+1425] + a; end
12'd1426: begin if(a[1426]==1) 
	 		intermediate[4095+1426:0+1426] <= intermediate[4095+1426:0+1426] + a; end
12'd1427: begin if(a[1427]==1) 
	 		intermediate[4095+1427:0+1427] <= intermediate[4095+1427:0+1427] + a; end
12'd1428: begin if(a[1428]==1) 
	 		intermediate[4095+1428:0+1428] <= intermediate[4095+1428:0+1428] + a; end
12'd1429: begin if(a[1429]==1) 
	 		intermediate[4095+1429:0+1429] <= intermediate[4095+1429:0+1429] + a; end
12'd1430: begin if(a[1430]==1) 
	 		intermediate[4095+1430:0+1430] <= intermediate[4095+1430:0+1430] + a; end
12'd1431: begin if(a[1431]==1) 
	 		intermediate[4095+1431:0+1431] <= intermediate[4095+1431:0+1431] + a; end
12'd1432: begin if(a[1432]==1) 
	 		intermediate[4095+1432:0+1432] <= intermediate[4095+1432:0+1432] + a; end
12'd1433: begin if(a[1433]==1) 
	 		intermediate[4095+1433:0+1433] <= intermediate[4095+1433:0+1433] + a; end
12'd1434: begin if(a[1434]==1) 
	 		intermediate[4095+1434:0+1434] <= intermediate[4095+1434:0+1434] + a; end
12'd1435: begin if(a[1435]==1) 
	 		intermediate[4095+1435:0+1435] <= intermediate[4095+1435:0+1435] + a; end
12'd1436: begin if(a[1436]==1) 
	 		intermediate[4095+1436:0+1436] <= intermediate[4095+1436:0+1436] + a; end
12'd1437: begin if(a[1437]==1) 
	 		intermediate[4095+1437:0+1437] <= intermediate[4095+1437:0+1437] + a; end
12'd1438: begin if(a[1438]==1) 
	 		intermediate[4095+1438:0+1438] <= intermediate[4095+1438:0+1438] + a; end
12'd1439: begin if(a[1439]==1) 
	 		intermediate[4095+1439:0+1439] <= intermediate[4095+1439:0+1439] + a; end
12'd1440: begin if(a[1440]==1) 
	 		intermediate[4095+1440:0+1440] <= intermediate[4095+1440:0+1440] + a; end
12'd1441: begin if(a[1441]==1) 
	 		intermediate[4095+1441:0+1441] <= intermediate[4095+1441:0+1441] + a; end
12'd1442: begin if(a[1442]==1) 
	 		intermediate[4095+1442:0+1442] <= intermediate[4095+1442:0+1442] + a; end
12'd1443: begin if(a[1443]==1) 
	 		intermediate[4095+1443:0+1443] <= intermediate[4095+1443:0+1443] + a; end
12'd1444: begin if(a[1444]==1) 
	 		intermediate[4095+1444:0+1444] <= intermediate[4095+1444:0+1444] + a; end
12'd1445: begin if(a[1445]==1) 
	 		intermediate[4095+1445:0+1445] <= intermediate[4095+1445:0+1445] + a; end
12'd1446: begin if(a[1446]==1) 
	 		intermediate[4095+1446:0+1446] <= intermediate[4095+1446:0+1446] + a; end
12'd1447: begin if(a[1447]==1) 
	 		intermediate[4095+1447:0+1447] <= intermediate[4095+1447:0+1447] + a; end
12'd1448: begin if(a[1448]==1) 
	 		intermediate[4095+1448:0+1448] <= intermediate[4095+1448:0+1448] + a; end
12'd1449: begin if(a[1449]==1) 
	 		intermediate[4095+1449:0+1449] <= intermediate[4095+1449:0+1449] + a; end
12'd1450: begin if(a[1450]==1) 
	 		intermediate[4095+1450:0+1450] <= intermediate[4095+1450:0+1450] + a; end
12'd1451: begin if(a[1451]==1) 
	 		intermediate[4095+1451:0+1451] <= intermediate[4095+1451:0+1451] + a; end
12'd1452: begin if(a[1452]==1) 
	 		intermediate[4095+1452:0+1452] <= intermediate[4095+1452:0+1452] + a; end
12'd1453: begin if(a[1453]==1) 
	 		intermediate[4095+1453:0+1453] <= intermediate[4095+1453:0+1453] + a; end
12'd1454: begin if(a[1454]==1) 
	 		intermediate[4095+1454:0+1454] <= intermediate[4095+1454:0+1454] + a; end
12'd1455: begin if(a[1455]==1) 
	 		intermediate[4095+1455:0+1455] <= intermediate[4095+1455:0+1455] + a; end
12'd1456: begin if(a[1456]==1) 
	 		intermediate[4095+1456:0+1456] <= intermediate[4095+1456:0+1456] + a; end
12'd1457: begin if(a[1457]==1) 
	 		intermediate[4095+1457:0+1457] <= intermediate[4095+1457:0+1457] + a; end
12'd1458: begin if(a[1458]==1) 
	 		intermediate[4095+1458:0+1458] <= intermediate[4095+1458:0+1458] + a; end
12'd1459: begin if(a[1459]==1) 
	 		intermediate[4095+1459:0+1459] <= intermediate[4095+1459:0+1459] + a; end
12'd1460: begin if(a[1460]==1) 
	 		intermediate[4095+1460:0+1460] <= intermediate[4095+1460:0+1460] + a; end
12'd1461: begin if(a[1461]==1) 
	 		intermediate[4095+1461:0+1461] <= intermediate[4095+1461:0+1461] + a; end
12'd1462: begin if(a[1462]==1) 
	 		intermediate[4095+1462:0+1462] <= intermediate[4095+1462:0+1462] + a; end
12'd1463: begin if(a[1463]==1) 
	 		intermediate[4095+1463:0+1463] <= intermediate[4095+1463:0+1463] + a; end
12'd1464: begin if(a[1464]==1) 
	 		intermediate[4095+1464:0+1464] <= intermediate[4095+1464:0+1464] + a; end
12'd1465: begin if(a[1465]==1) 
	 		intermediate[4095+1465:0+1465] <= intermediate[4095+1465:0+1465] + a; end
12'd1466: begin if(a[1466]==1) 
	 		intermediate[4095+1466:0+1466] <= intermediate[4095+1466:0+1466] + a; end
12'd1467: begin if(a[1467]==1) 
	 		intermediate[4095+1467:0+1467] <= intermediate[4095+1467:0+1467] + a; end
12'd1468: begin if(a[1468]==1) 
	 		intermediate[4095+1468:0+1468] <= intermediate[4095+1468:0+1468] + a; end
12'd1469: begin if(a[1469]==1) 
	 		intermediate[4095+1469:0+1469] <= intermediate[4095+1469:0+1469] + a; end
12'd1470: begin if(a[1470]==1) 
	 		intermediate[4095+1470:0+1470] <= intermediate[4095+1470:0+1470] + a; end
12'd1471: begin if(a[1471]==1) 
	 		intermediate[4095+1471:0+1471] <= intermediate[4095+1471:0+1471] + a; end
12'd1472: begin if(a[1472]==1) 
	 		intermediate[4095+1472:0+1472] <= intermediate[4095+1472:0+1472] + a; end
12'd1473: begin if(a[1473]==1) 
	 		intermediate[4095+1473:0+1473] <= intermediate[4095+1473:0+1473] + a; end
12'd1474: begin if(a[1474]==1) 
	 		intermediate[4095+1474:0+1474] <= intermediate[4095+1474:0+1474] + a; end
12'd1475: begin if(a[1475]==1) 
	 		intermediate[4095+1475:0+1475] <= intermediate[4095+1475:0+1475] + a; end
12'd1476: begin if(a[1476]==1) 
	 		intermediate[4095+1476:0+1476] <= intermediate[4095+1476:0+1476] + a; end
12'd1477: begin if(a[1477]==1) 
	 		intermediate[4095+1477:0+1477] <= intermediate[4095+1477:0+1477] + a; end
12'd1478: begin if(a[1478]==1) 
	 		intermediate[4095+1478:0+1478] <= intermediate[4095+1478:0+1478] + a; end
12'd1479: begin if(a[1479]==1) 
	 		intermediate[4095+1479:0+1479] <= intermediate[4095+1479:0+1479] + a; end
12'd1480: begin if(a[1480]==1) 
	 		intermediate[4095+1480:0+1480] <= intermediate[4095+1480:0+1480] + a; end
12'd1481: begin if(a[1481]==1) 
	 		intermediate[4095+1481:0+1481] <= intermediate[4095+1481:0+1481] + a; end
12'd1482: begin if(a[1482]==1) 
	 		intermediate[4095+1482:0+1482] <= intermediate[4095+1482:0+1482] + a; end
12'd1483: begin if(a[1483]==1) 
	 		intermediate[4095+1483:0+1483] <= intermediate[4095+1483:0+1483] + a; end
12'd1484: begin if(a[1484]==1) 
	 		intermediate[4095+1484:0+1484] <= intermediate[4095+1484:0+1484] + a; end
12'd1485: begin if(a[1485]==1) 
	 		intermediate[4095+1485:0+1485] <= intermediate[4095+1485:0+1485] + a; end
12'd1486: begin if(a[1486]==1) 
	 		intermediate[4095+1486:0+1486] <= intermediate[4095+1486:0+1486] + a; end
12'd1487: begin if(a[1487]==1) 
	 		intermediate[4095+1487:0+1487] <= intermediate[4095+1487:0+1487] + a; end
12'd1488: begin if(a[1488]==1) 
	 		intermediate[4095+1488:0+1488] <= intermediate[4095+1488:0+1488] + a; end
12'd1489: begin if(a[1489]==1) 
	 		intermediate[4095+1489:0+1489] <= intermediate[4095+1489:0+1489] + a; end
12'd1490: begin if(a[1490]==1) 
	 		intermediate[4095+1490:0+1490] <= intermediate[4095+1490:0+1490] + a; end
12'd1491: begin if(a[1491]==1) 
	 		intermediate[4095+1491:0+1491] <= intermediate[4095+1491:0+1491] + a; end
12'd1492: begin if(a[1492]==1) 
	 		intermediate[4095+1492:0+1492] <= intermediate[4095+1492:0+1492] + a; end
12'd1493: begin if(a[1493]==1) 
	 		intermediate[4095+1493:0+1493] <= intermediate[4095+1493:0+1493] + a; end
12'd1494: begin if(a[1494]==1) 
	 		intermediate[4095+1494:0+1494] <= intermediate[4095+1494:0+1494] + a; end
12'd1495: begin if(a[1495]==1) 
	 		intermediate[4095+1495:0+1495] <= intermediate[4095+1495:0+1495] + a; end
12'd1496: begin if(a[1496]==1) 
	 		intermediate[4095+1496:0+1496] <= intermediate[4095+1496:0+1496] + a; end
12'd1497: begin if(a[1497]==1) 
	 		intermediate[4095+1497:0+1497] <= intermediate[4095+1497:0+1497] + a; end
12'd1498: begin if(a[1498]==1) 
	 		intermediate[4095+1498:0+1498] <= intermediate[4095+1498:0+1498] + a; end
12'd1499: begin if(a[1499]==1) 
	 		intermediate[4095+1499:0+1499] <= intermediate[4095+1499:0+1499] + a; end
12'd1500: begin if(a[1500]==1) 
	 		intermediate[4095+1500:0+1500] <= intermediate[4095+1500:0+1500] + a; end
12'd1501: begin if(a[1501]==1) 
	 		intermediate[4095+1501:0+1501] <= intermediate[4095+1501:0+1501] + a; end
12'd1502: begin if(a[1502]==1) 
	 		intermediate[4095+1502:0+1502] <= intermediate[4095+1502:0+1502] + a; end
12'd1503: begin if(a[1503]==1) 
	 		intermediate[4095+1503:0+1503] <= intermediate[4095+1503:0+1503] + a; end
12'd1504: begin if(a[1504]==1) 
	 		intermediate[4095+1504:0+1504] <= intermediate[4095+1504:0+1504] + a; end
12'd1505: begin if(a[1505]==1) 
	 		intermediate[4095+1505:0+1505] <= intermediate[4095+1505:0+1505] + a; end
12'd1506: begin if(a[1506]==1) 
	 		intermediate[4095+1506:0+1506] <= intermediate[4095+1506:0+1506] + a; end
12'd1507: begin if(a[1507]==1) 
	 		intermediate[4095+1507:0+1507] <= intermediate[4095+1507:0+1507] + a; end
12'd1508: begin if(a[1508]==1) 
	 		intermediate[4095+1508:0+1508] <= intermediate[4095+1508:0+1508] + a; end
12'd1509: begin if(a[1509]==1) 
	 		intermediate[4095+1509:0+1509] <= intermediate[4095+1509:0+1509] + a; end
12'd1510: begin if(a[1510]==1) 
	 		intermediate[4095+1510:0+1510] <= intermediate[4095+1510:0+1510] + a; end
12'd1511: begin if(a[1511]==1) 
	 		intermediate[4095+1511:0+1511] <= intermediate[4095+1511:0+1511] + a; end
12'd1512: begin if(a[1512]==1) 
	 		intermediate[4095+1512:0+1512] <= intermediate[4095+1512:0+1512] + a; end
12'd1513: begin if(a[1513]==1) 
	 		intermediate[4095+1513:0+1513] <= intermediate[4095+1513:0+1513] + a; end
12'd1514: begin if(a[1514]==1) 
	 		intermediate[4095+1514:0+1514] <= intermediate[4095+1514:0+1514] + a; end
12'd1515: begin if(a[1515]==1) 
	 		intermediate[4095+1515:0+1515] <= intermediate[4095+1515:0+1515] + a; end
12'd1516: begin if(a[1516]==1) 
	 		intermediate[4095+1516:0+1516] <= intermediate[4095+1516:0+1516] + a; end
12'd1517: begin if(a[1517]==1) 
	 		intermediate[4095+1517:0+1517] <= intermediate[4095+1517:0+1517] + a; end
12'd1518: begin if(a[1518]==1) 
	 		intermediate[4095+1518:0+1518] <= intermediate[4095+1518:0+1518] + a; end
12'd1519: begin if(a[1519]==1) 
	 		intermediate[4095+1519:0+1519] <= intermediate[4095+1519:0+1519] + a; end
12'd1520: begin if(a[1520]==1) 
	 		intermediate[4095+1520:0+1520] <= intermediate[4095+1520:0+1520] + a; end
12'd1521: begin if(a[1521]==1) 
	 		intermediate[4095+1521:0+1521] <= intermediate[4095+1521:0+1521] + a; end
12'd1522: begin if(a[1522]==1) 
	 		intermediate[4095+1522:0+1522] <= intermediate[4095+1522:0+1522] + a; end
12'd1523: begin if(a[1523]==1) 
	 		intermediate[4095+1523:0+1523] <= intermediate[4095+1523:0+1523] + a; end
12'd1524: begin if(a[1524]==1) 
	 		intermediate[4095+1524:0+1524] <= intermediate[4095+1524:0+1524] + a; end
12'd1525: begin if(a[1525]==1) 
	 		intermediate[4095+1525:0+1525] <= intermediate[4095+1525:0+1525] + a; end
12'd1526: begin if(a[1526]==1) 
	 		intermediate[4095+1526:0+1526] <= intermediate[4095+1526:0+1526] + a; end
12'd1527: begin if(a[1527]==1) 
	 		intermediate[4095+1527:0+1527] <= intermediate[4095+1527:0+1527] + a; end
12'd1528: begin if(a[1528]==1) 
	 		intermediate[4095+1528:0+1528] <= intermediate[4095+1528:0+1528] + a; end
12'd1529: begin if(a[1529]==1) 
	 		intermediate[4095+1529:0+1529] <= intermediate[4095+1529:0+1529] + a; end
12'd1530: begin if(a[1530]==1) 
	 		intermediate[4095+1530:0+1530] <= intermediate[4095+1530:0+1530] + a; end
12'd1531: begin if(a[1531]==1) 
	 		intermediate[4095+1531:0+1531] <= intermediate[4095+1531:0+1531] + a; end
12'd1532: begin if(a[1532]==1) 
	 		intermediate[4095+1532:0+1532] <= intermediate[4095+1532:0+1532] + a; end
12'd1533: begin if(a[1533]==1) 
	 		intermediate[4095+1533:0+1533] <= intermediate[4095+1533:0+1533] + a; end
12'd1534: begin if(a[1534]==1) 
	 		intermediate[4095+1534:0+1534] <= intermediate[4095+1534:0+1534] + a; end
12'd1535: begin if(a[1535]==1) 
	 		intermediate[4095+1535:0+1535] <= intermediate[4095+1535:0+1535] + a; end
12'd1536: begin if(a[1536]==1) 
	 		intermediate[4095+1536:0+1536] <= intermediate[4095+1536:0+1536] + a; end
12'd1537: begin if(a[1537]==1) 
	 		intermediate[4095+1537:0+1537] <= intermediate[4095+1537:0+1537] + a; end
12'd1538: begin if(a[1538]==1) 
	 		intermediate[4095+1538:0+1538] <= intermediate[4095+1538:0+1538] + a; end
12'd1539: begin if(a[1539]==1) 
	 		intermediate[4095+1539:0+1539] <= intermediate[4095+1539:0+1539] + a; end
12'd1540: begin if(a[1540]==1) 
	 		intermediate[4095+1540:0+1540] <= intermediate[4095+1540:0+1540] + a; end
12'd1541: begin if(a[1541]==1) 
	 		intermediate[4095+1541:0+1541] <= intermediate[4095+1541:0+1541] + a; end
12'd1542: begin if(a[1542]==1) 
	 		intermediate[4095+1542:0+1542] <= intermediate[4095+1542:0+1542] + a; end
12'd1543: begin if(a[1543]==1) 
	 		intermediate[4095+1543:0+1543] <= intermediate[4095+1543:0+1543] + a; end
12'd1544: begin if(a[1544]==1) 
	 		intermediate[4095+1544:0+1544] <= intermediate[4095+1544:0+1544] + a; end
12'd1545: begin if(a[1545]==1) 
	 		intermediate[4095+1545:0+1545] <= intermediate[4095+1545:0+1545] + a; end
12'd1546: begin if(a[1546]==1) 
	 		intermediate[4095+1546:0+1546] <= intermediate[4095+1546:0+1546] + a; end
12'd1547: begin if(a[1547]==1) 
	 		intermediate[4095+1547:0+1547] <= intermediate[4095+1547:0+1547] + a; end
12'd1548: begin if(a[1548]==1) 
	 		intermediate[4095+1548:0+1548] <= intermediate[4095+1548:0+1548] + a; end
12'd1549: begin if(a[1549]==1) 
	 		intermediate[4095+1549:0+1549] <= intermediate[4095+1549:0+1549] + a; end
12'd1550: begin if(a[1550]==1) 
	 		intermediate[4095+1550:0+1550] <= intermediate[4095+1550:0+1550] + a; end
12'd1551: begin if(a[1551]==1) 
	 		intermediate[4095+1551:0+1551] <= intermediate[4095+1551:0+1551] + a; end
12'd1552: begin if(a[1552]==1) 
	 		intermediate[4095+1552:0+1552] <= intermediate[4095+1552:0+1552] + a; end
12'd1553: begin if(a[1553]==1) 
	 		intermediate[4095+1553:0+1553] <= intermediate[4095+1553:0+1553] + a; end
12'd1554: begin if(a[1554]==1) 
	 		intermediate[4095+1554:0+1554] <= intermediate[4095+1554:0+1554] + a; end
12'd1555: begin if(a[1555]==1) 
	 		intermediate[4095+1555:0+1555] <= intermediate[4095+1555:0+1555] + a; end
12'd1556: begin if(a[1556]==1) 
	 		intermediate[4095+1556:0+1556] <= intermediate[4095+1556:0+1556] + a; end
12'd1557: begin if(a[1557]==1) 
	 		intermediate[4095+1557:0+1557] <= intermediate[4095+1557:0+1557] + a; end
12'd1558: begin if(a[1558]==1) 
	 		intermediate[4095+1558:0+1558] <= intermediate[4095+1558:0+1558] + a; end
12'd1559: begin if(a[1559]==1) 
	 		intermediate[4095+1559:0+1559] <= intermediate[4095+1559:0+1559] + a; end
12'd1560: begin if(a[1560]==1) 
	 		intermediate[4095+1560:0+1560] <= intermediate[4095+1560:0+1560] + a; end
12'd1561: begin if(a[1561]==1) 
	 		intermediate[4095+1561:0+1561] <= intermediate[4095+1561:0+1561] + a; end
12'd1562: begin if(a[1562]==1) 
	 		intermediate[4095+1562:0+1562] <= intermediate[4095+1562:0+1562] + a; end
12'd1563: begin if(a[1563]==1) 
	 		intermediate[4095+1563:0+1563] <= intermediate[4095+1563:0+1563] + a; end
12'd1564: begin if(a[1564]==1) 
	 		intermediate[4095+1564:0+1564] <= intermediate[4095+1564:0+1564] + a; end
12'd1565: begin if(a[1565]==1) 
	 		intermediate[4095+1565:0+1565] <= intermediate[4095+1565:0+1565] + a; end
12'd1566: begin if(a[1566]==1) 
	 		intermediate[4095+1566:0+1566] <= intermediate[4095+1566:0+1566] + a; end
12'd1567: begin if(a[1567]==1) 
	 		intermediate[4095+1567:0+1567] <= intermediate[4095+1567:0+1567] + a; end
12'd1568: begin if(a[1568]==1) 
	 		intermediate[4095+1568:0+1568] <= intermediate[4095+1568:0+1568] + a; end
12'd1569: begin if(a[1569]==1) 
	 		intermediate[4095+1569:0+1569] <= intermediate[4095+1569:0+1569] + a; end
12'd1570: begin if(a[1570]==1) 
	 		intermediate[4095+1570:0+1570] <= intermediate[4095+1570:0+1570] + a; end
12'd1571: begin if(a[1571]==1) 
	 		intermediate[4095+1571:0+1571] <= intermediate[4095+1571:0+1571] + a; end
12'd1572: begin if(a[1572]==1) 
	 		intermediate[4095+1572:0+1572] <= intermediate[4095+1572:0+1572] + a; end
12'd1573: begin if(a[1573]==1) 
	 		intermediate[4095+1573:0+1573] <= intermediate[4095+1573:0+1573] + a; end
12'd1574: begin if(a[1574]==1) 
	 		intermediate[4095+1574:0+1574] <= intermediate[4095+1574:0+1574] + a; end
12'd1575: begin if(a[1575]==1) 
	 		intermediate[4095+1575:0+1575] <= intermediate[4095+1575:0+1575] + a; end
12'd1576: begin if(a[1576]==1) 
	 		intermediate[4095+1576:0+1576] <= intermediate[4095+1576:0+1576] + a; end
12'd1577: begin if(a[1577]==1) 
	 		intermediate[4095+1577:0+1577] <= intermediate[4095+1577:0+1577] + a; end
12'd1578: begin if(a[1578]==1) 
	 		intermediate[4095+1578:0+1578] <= intermediate[4095+1578:0+1578] + a; end
12'd1579: begin if(a[1579]==1) 
	 		intermediate[4095+1579:0+1579] <= intermediate[4095+1579:0+1579] + a; end
12'd1580: begin if(a[1580]==1) 
	 		intermediate[4095+1580:0+1580] <= intermediate[4095+1580:0+1580] + a; end
12'd1581: begin if(a[1581]==1) 
	 		intermediate[4095+1581:0+1581] <= intermediate[4095+1581:0+1581] + a; end
12'd1582: begin if(a[1582]==1) 
	 		intermediate[4095+1582:0+1582] <= intermediate[4095+1582:0+1582] + a; end
12'd1583: begin if(a[1583]==1) 
	 		intermediate[4095+1583:0+1583] <= intermediate[4095+1583:0+1583] + a; end
12'd1584: begin if(a[1584]==1) 
	 		intermediate[4095+1584:0+1584] <= intermediate[4095+1584:0+1584] + a; end
12'd1585: begin if(a[1585]==1) 
	 		intermediate[4095+1585:0+1585] <= intermediate[4095+1585:0+1585] + a; end
12'd1586: begin if(a[1586]==1) 
	 		intermediate[4095+1586:0+1586] <= intermediate[4095+1586:0+1586] + a; end
12'd1587: begin if(a[1587]==1) 
	 		intermediate[4095+1587:0+1587] <= intermediate[4095+1587:0+1587] + a; end
12'd1588: begin if(a[1588]==1) 
	 		intermediate[4095+1588:0+1588] <= intermediate[4095+1588:0+1588] + a; end
12'd1589: begin if(a[1589]==1) 
	 		intermediate[4095+1589:0+1589] <= intermediate[4095+1589:0+1589] + a; end
12'd1590: begin if(a[1590]==1) 
	 		intermediate[4095+1590:0+1590] <= intermediate[4095+1590:0+1590] + a; end
12'd1591: begin if(a[1591]==1) 
	 		intermediate[4095+1591:0+1591] <= intermediate[4095+1591:0+1591] + a; end
12'd1592: begin if(a[1592]==1) 
	 		intermediate[4095+1592:0+1592] <= intermediate[4095+1592:0+1592] + a; end
12'd1593: begin if(a[1593]==1) 
	 		intermediate[4095+1593:0+1593] <= intermediate[4095+1593:0+1593] + a; end
12'd1594: begin if(a[1594]==1) 
	 		intermediate[4095+1594:0+1594] <= intermediate[4095+1594:0+1594] + a; end
12'd1595: begin if(a[1595]==1) 
	 		intermediate[4095+1595:0+1595] <= intermediate[4095+1595:0+1595] + a; end
12'd1596: begin if(a[1596]==1) 
	 		intermediate[4095+1596:0+1596] <= intermediate[4095+1596:0+1596] + a; end
12'd1597: begin if(a[1597]==1) 
	 		intermediate[4095+1597:0+1597] <= intermediate[4095+1597:0+1597] + a; end
12'd1598: begin if(a[1598]==1) 
	 		intermediate[4095+1598:0+1598] <= intermediate[4095+1598:0+1598] + a; end
12'd1599: begin if(a[1599]==1) 
	 		intermediate[4095+1599:0+1599] <= intermediate[4095+1599:0+1599] + a; end
12'd1600: begin if(a[1600]==1) 
	 		intermediate[4095+1600:0+1600] <= intermediate[4095+1600:0+1600] + a; end
12'd1601: begin if(a[1601]==1) 
	 		intermediate[4095+1601:0+1601] <= intermediate[4095+1601:0+1601] + a; end
12'd1602: begin if(a[1602]==1) 
	 		intermediate[4095+1602:0+1602] <= intermediate[4095+1602:0+1602] + a; end
12'd1603: begin if(a[1603]==1) 
	 		intermediate[4095+1603:0+1603] <= intermediate[4095+1603:0+1603] + a; end
12'd1604: begin if(a[1604]==1) 
	 		intermediate[4095+1604:0+1604] <= intermediate[4095+1604:0+1604] + a; end
12'd1605: begin if(a[1605]==1) 
	 		intermediate[4095+1605:0+1605] <= intermediate[4095+1605:0+1605] + a; end
12'd1606: begin if(a[1606]==1) 
	 		intermediate[4095+1606:0+1606] <= intermediate[4095+1606:0+1606] + a; end
12'd1607: begin if(a[1607]==1) 
	 		intermediate[4095+1607:0+1607] <= intermediate[4095+1607:0+1607] + a; end
12'd1608: begin if(a[1608]==1) 
	 		intermediate[4095+1608:0+1608] <= intermediate[4095+1608:0+1608] + a; end
12'd1609: begin if(a[1609]==1) 
	 		intermediate[4095+1609:0+1609] <= intermediate[4095+1609:0+1609] + a; end
12'd1610: begin if(a[1610]==1) 
	 		intermediate[4095+1610:0+1610] <= intermediate[4095+1610:0+1610] + a; end
12'd1611: begin if(a[1611]==1) 
	 		intermediate[4095+1611:0+1611] <= intermediate[4095+1611:0+1611] + a; end
12'd1612: begin if(a[1612]==1) 
	 		intermediate[4095+1612:0+1612] <= intermediate[4095+1612:0+1612] + a; end
12'd1613: begin if(a[1613]==1) 
	 		intermediate[4095+1613:0+1613] <= intermediate[4095+1613:0+1613] + a; end
12'd1614: begin if(a[1614]==1) 
	 		intermediate[4095+1614:0+1614] <= intermediate[4095+1614:0+1614] + a; end
12'd1615: begin if(a[1615]==1) 
	 		intermediate[4095+1615:0+1615] <= intermediate[4095+1615:0+1615] + a; end
12'd1616: begin if(a[1616]==1) 
	 		intermediate[4095+1616:0+1616] <= intermediate[4095+1616:0+1616] + a; end
12'd1617: begin if(a[1617]==1) 
	 		intermediate[4095+1617:0+1617] <= intermediate[4095+1617:0+1617] + a; end
12'd1618: begin if(a[1618]==1) 
	 		intermediate[4095+1618:0+1618] <= intermediate[4095+1618:0+1618] + a; end
12'd1619: begin if(a[1619]==1) 
	 		intermediate[4095+1619:0+1619] <= intermediate[4095+1619:0+1619] + a; end
12'd1620: begin if(a[1620]==1) 
	 		intermediate[4095+1620:0+1620] <= intermediate[4095+1620:0+1620] + a; end
12'd1621: begin if(a[1621]==1) 
	 		intermediate[4095+1621:0+1621] <= intermediate[4095+1621:0+1621] + a; end
12'd1622: begin if(a[1622]==1) 
	 		intermediate[4095+1622:0+1622] <= intermediate[4095+1622:0+1622] + a; end
12'd1623: begin if(a[1623]==1) 
	 		intermediate[4095+1623:0+1623] <= intermediate[4095+1623:0+1623] + a; end
12'd1624: begin if(a[1624]==1) 
	 		intermediate[4095+1624:0+1624] <= intermediate[4095+1624:0+1624] + a; end
12'd1625: begin if(a[1625]==1) 
	 		intermediate[4095+1625:0+1625] <= intermediate[4095+1625:0+1625] + a; end
12'd1626: begin if(a[1626]==1) 
	 		intermediate[4095+1626:0+1626] <= intermediate[4095+1626:0+1626] + a; end
12'd1627: begin if(a[1627]==1) 
	 		intermediate[4095+1627:0+1627] <= intermediate[4095+1627:0+1627] + a; end
12'd1628: begin if(a[1628]==1) 
	 		intermediate[4095+1628:0+1628] <= intermediate[4095+1628:0+1628] + a; end
12'd1629: begin if(a[1629]==1) 
	 		intermediate[4095+1629:0+1629] <= intermediate[4095+1629:0+1629] + a; end
12'd1630: begin if(a[1630]==1) 
	 		intermediate[4095+1630:0+1630] <= intermediate[4095+1630:0+1630] + a; end
12'd1631: begin if(a[1631]==1) 
	 		intermediate[4095+1631:0+1631] <= intermediate[4095+1631:0+1631] + a; end
12'd1632: begin if(a[1632]==1) 
	 		intermediate[4095+1632:0+1632] <= intermediate[4095+1632:0+1632] + a; end
12'd1633: begin if(a[1633]==1) 
	 		intermediate[4095+1633:0+1633] <= intermediate[4095+1633:0+1633] + a; end
12'd1634: begin if(a[1634]==1) 
	 		intermediate[4095+1634:0+1634] <= intermediate[4095+1634:0+1634] + a; end
12'd1635: begin if(a[1635]==1) 
	 		intermediate[4095+1635:0+1635] <= intermediate[4095+1635:0+1635] + a; end
12'd1636: begin if(a[1636]==1) 
	 		intermediate[4095+1636:0+1636] <= intermediate[4095+1636:0+1636] + a; end
12'd1637: begin if(a[1637]==1) 
	 		intermediate[4095+1637:0+1637] <= intermediate[4095+1637:0+1637] + a; end
12'd1638: begin if(a[1638]==1) 
	 		intermediate[4095+1638:0+1638] <= intermediate[4095+1638:0+1638] + a; end
12'd1639: begin if(a[1639]==1) 
	 		intermediate[4095+1639:0+1639] <= intermediate[4095+1639:0+1639] + a; end
12'd1640: begin if(a[1640]==1) 
	 		intermediate[4095+1640:0+1640] <= intermediate[4095+1640:0+1640] + a; end
12'd1641: begin if(a[1641]==1) 
	 		intermediate[4095+1641:0+1641] <= intermediate[4095+1641:0+1641] + a; end
12'd1642: begin if(a[1642]==1) 
	 		intermediate[4095+1642:0+1642] <= intermediate[4095+1642:0+1642] + a; end
12'd1643: begin if(a[1643]==1) 
	 		intermediate[4095+1643:0+1643] <= intermediate[4095+1643:0+1643] + a; end
12'd1644: begin if(a[1644]==1) 
	 		intermediate[4095+1644:0+1644] <= intermediate[4095+1644:0+1644] + a; end
12'd1645: begin if(a[1645]==1) 
	 		intermediate[4095+1645:0+1645] <= intermediate[4095+1645:0+1645] + a; end
12'd1646: begin if(a[1646]==1) 
	 		intermediate[4095+1646:0+1646] <= intermediate[4095+1646:0+1646] + a; end
12'd1647: begin if(a[1647]==1) 
	 		intermediate[4095+1647:0+1647] <= intermediate[4095+1647:0+1647] + a; end
12'd1648: begin if(a[1648]==1) 
	 		intermediate[4095+1648:0+1648] <= intermediate[4095+1648:0+1648] + a; end
12'd1649: begin if(a[1649]==1) 
	 		intermediate[4095+1649:0+1649] <= intermediate[4095+1649:0+1649] + a; end
12'd1650: begin if(a[1650]==1) 
	 		intermediate[4095+1650:0+1650] <= intermediate[4095+1650:0+1650] + a; end
12'd1651: begin if(a[1651]==1) 
	 		intermediate[4095+1651:0+1651] <= intermediate[4095+1651:0+1651] + a; end
12'd1652: begin if(a[1652]==1) 
	 		intermediate[4095+1652:0+1652] <= intermediate[4095+1652:0+1652] + a; end
12'd1653: begin if(a[1653]==1) 
	 		intermediate[4095+1653:0+1653] <= intermediate[4095+1653:0+1653] + a; end
12'd1654: begin if(a[1654]==1) 
	 		intermediate[4095+1654:0+1654] <= intermediate[4095+1654:0+1654] + a; end
12'd1655: begin if(a[1655]==1) 
	 		intermediate[4095+1655:0+1655] <= intermediate[4095+1655:0+1655] + a; end
12'd1656: begin if(a[1656]==1) 
	 		intermediate[4095+1656:0+1656] <= intermediate[4095+1656:0+1656] + a; end
12'd1657: begin if(a[1657]==1) 
	 		intermediate[4095+1657:0+1657] <= intermediate[4095+1657:0+1657] + a; end
12'd1658: begin if(a[1658]==1) 
	 		intermediate[4095+1658:0+1658] <= intermediate[4095+1658:0+1658] + a; end
12'd1659: begin if(a[1659]==1) 
	 		intermediate[4095+1659:0+1659] <= intermediate[4095+1659:0+1659] + a; end
12'd1660: begin if(a[1660]==1) 
	 		intermediate[4095+1660:0+1660] <= intermediate[4095+1660:0+1660] + a; end
12'd1661: begin if(a[1661]==1) 
	 		intermediate[4095+1661:0+1661] <= intermediate[4095+1661:0+1661] + a; end
12'd1662: begin if(a[1662]==1) 
	 		intermediate[4095+1662:0+1662] <= intermediate[4095+1662:0+1662] + a; end
12'd1663: begin if(a[1663]==1) 
	 		intermediate[4095+1663:0+1663] <= intermediate[4095+1663:0+1663] + a; end
12'd1664: begin if(a[1664]==1) 
	 		intermediate[4095+1664:0+1664] <= intermediate[4095+1664:0+1664] + a; end
12'd1665: begin if(a[1665]==1) 
	 		intermediate[4095+1665:0+1665] <= intermediate[4095+1665:0+1665] + a; end
12'd1666: begin if(a[1666]==1) 
	 		intermediate[4095+1666:0+1666] <= intermediate[4095+1666:0+1666] + a; end
12'd1667: begin if(a[1667]==1) 
	 		intermediate[4095+1667:0+1667] <= intermediate[4095+1667:0+1667] + a; end
12'd1668: begin if(a[1668]==1) 
	 		intermediate[4095+1668:0+1668] <= intermediate[4095+1668:0+1668] + a; end
12'd1669: begin if(a[1669]==1) 
	 		intermediate[4095+1669:0+1669] <= intermediate[4095+1669:0+1669] + a; end
12'd1670: begin if(a[1670]==1) 
	 		intermediate[4095+1670:0+1670] <= intermediate[4095+1670:0+1670] + a; end
12'd1671: begin if(a[1671]==1) 
	 		intermediate[4095+1671:0+1671] <= intermediate[4095+1671:0+1671] + a; end
12'd1672: begin if(a[1672]==1) 
	 		intermediate[4095+1672:0+1672] <= intermediate[4095+1672:0+1672] + a; end
12'd1673: begin if(a[1673]==1) 
	 		intermediate[4095+1673:0+1673] <= intermediate[4095+1673:0+1673] + a; end
12'd1674: begin if(a[1674]==1) 
	 		intermediate[4095+1674:0+1674] <= intermediate[4095+1674:0+1674] + a; end
12'd1675: begin if(a[1675]==1) 
	 		intermediate[4095+1675:0+1675] <= intermediate[4095+1675:0+1675] + a; end
12'd1676: begin if(a[1676]==1) 
	 		intermediate[4095+1676:0+1676] <= intermediate[4095+1676:0+1676] + a; end
12'd1677: begin if(a[1677]==1) 
	 		intermediate[4095+1677:0+1677] <= intermediate[4095+1677:0+1677] + a; end
12'd1678: begin if(a[1678]==1) 
	 		intermediate[4095+1678:0+1678] <= intermediate[4095+1678:0+1678] + a; end
12'd1679: begin if(a[1679]==1) 
	 		intermediate[4095+1679:0+1679] <= intermediate[4095+1679:0+1679] + a; end
12'd1680: begin if(a[1680]==1) 
	 		intermediate[4095+1680:0+1680] <= intermediate[4095+1680:0+1680] + a; end
12'd1681: begin if(a[1681]==1) 
	 		intermediate[4095+1681:0+1681] <= intermediate[4095+1681:0+1681] + a; end
12'd1682: begin if(a[1682]==1) 
	 		intermediate[4095+1682:0+1682] <= intermediate[4095+1682:0+1682] + a; end
12'd1683: begin if(a[1683]==1) 
	 		intermediate[4095+1683:0+1683] <= intermediate[4095+1683:0+1683] + a; end
12'd1684: begin if(a[1684]==1) 
	 		intermediate[4095+1684:0+1684] <= intermediate[4095+1684:0+1684] + a; end
12'd1685: begin if(a[1685]==1) 
	 		intermediate[4095+1685:0+1685] <= intermediate[4095+1685:0+1685] + a; end
12'd1686: begin if(a[1686]==1) 
	 		intermediate[4095+1686:0+1686] <= intermediate[4095+1686:0+1686] + a; end
12'd1687: begin if(a[1687]==1) 
	 		intermediate[4095+1687:0+1687] <= intermediate[4095+1687:0+1687] + a; end
12'd1688: begin if(a[1688]==1) 
	 		intermediate[4095+1688:0+1688] <= intermediate[4095+1688:0+1688] + a; end
12'd1689: begin if(a[1689]==1) 
	 		intermediate[4095+1689:0+1689] <= intermediate[4095+1689:0+1689] + a; end
12'd1690: begin if(a[1690]==1) 
	 		intermediate[4095+1690:0+1690] <= intermediate[4095+1690:0+1690] + a; end
12'd1691: begin if(a[1691]==1) 
	 		intermediate[4095+1691:0+1691] <= intermediate[4095+1691:0+1691] + a; end
12'd1692: begin if(a[1692]==1) 
	 		intermediate[4095+1692:0+1692] <= intermediate[4095+1692:0+1692] + a; end
12'd1693: begin if(a[1693]==1) 
	 		intermediate[4095+1693:0+1693] <= intermediate[4095+1693:0+1693] + a; end
12'd1694: begin if(a[1694]==1) 
	 		intermediate[4095+1694:0+1694] <= intermediate[4095+1694:0+1694] + a; end
12'd1695: begin if(a[1695]==1) 
	 		intermediate[4095+1695:0+1695] <= intermediate[4095+1695:0+1695] + a; end
12'd1696: begin if(a[1696]==1) 
	 		intermediate[4095+1696:0+1696] <= intermediate[4095+1696:0+1696] + a; end
12'd1697: begin if(a[1697]==1) 
	 		intermediate[4095+1697:0+1697] <= intermediate[4095+1697:0+1697] + a; end
12'd1698: begin if(a[1698]==1) 
	 		intermediate[4095+1698:0+1698] <= intermediate[4095+1698:0+1698] + a; end
12'd1699: begin if(a[1699]==1) 
	 		intermediate[4095+1699:0+1699] <= intermediate[4095+1699:0+1699] + a; end
12'd1700: begin if(a[1700]==1) 
	 		intermediate[4095+1700:0+1700] <= intermediate[4095+1700:0+1700] + a; end
12'd1701: begin if(a[1701]==1) 
	 		intermediate[4095+1701:0+1701] <= intermediate[4095+1701:0+1701] + a; end
12'd1702: begin if(a[1702]==1) 
	 		intermediate[4095+1702:0+1702] <= intermediate[4095+1702:0+1702] + a; end
12'd1703: begin if(a[1703]==1) 
	 		intermediate[4095+1703:0+1703] <= intermediate[4095+1703:0+1703] + a; end
12'd1704: begin if(a[1704]==1) 
	 		intermediate[4095+1704:0+1704] <= intermediate[4095+1704:0+1704] + a; end
12'd1705: begin if(a[1705]==1) 
	 		intermediate[4095+1705:0+1705] <= intermediate[4095+1705:0+1705] + a; end
12'd1706: begin if(a[1706]==1) 
	 		intermediate[4095+1706:0+1706] <= intermediate[4095+1706:0+1706] + a; end
12'd1707: begin if(a[1707]==1) 
	 		intermediate[4095+1707:0+1707] <= intermediate[4095+1707:0+1707] + a; end
12'd1708: begin if(a[1708]==1) 
	 		intermediate[4095+1708:0+1708] <= intermediate[4095+1708:0+1708] + a; end
12'd1709: begin if(a[1709]==1) 
	 		intermediate[4095+1709:0+1709] <= intermediate[4095+1709:0+1709] + a; end
12'd1710: begin if(a[1710]==1) 
	 		intermediate[4095+1710:0+1710] <= intermediate[4095+1710:0+1710] + a; end
12'd1711: begin if(a[1711]==1) 
	 		intermediate[4095+1711:0+1711] <= intermediate[4095+1711:0+1711] + a; end
12'd1712: begin if(a[1712]==1) 
	 		intermediate[4095+1712:0+1712] <= intermediate[4095+1712:0+1712] + a; end
12'd1713: begin if(a[1713]==1) 
	 		intermediate[4095+1713:0+1713] <= intermediate[4095+1713:0+1713] + a; end
12'd1714: begin if(a[1714]==1) 
	 		intermediate[4095+1714:0+1714] <= intermediate[4095+1714:0+1714] + a; end
12'd1715: begin if(a[1715]==1) 
	 		intermediate[4095+1715:0+1715] <= intermediate[4095+1715:0+1715] + a; end
12'd1716: begin if(a[1716]==1) 
	 		intermediate[4095+1716:0+1716] <= intermediate[4095+1716:0+1716] + a; end
12'd1717: begin if(a[1717]==1) 
	 		intermediate[4095+1717:0+1717] <= intermediate[4095+1717:0+1717] + a; end
12'd1718: begin if(a[1718]==1) 
	 		intermediate[4095+1718:0+1718] <= intermediate[4095+1718:0+1718] + a; end
12'd1719: begin if(a[1719]==1) 
	 		intermediate[4095+1719:0+1719] <= intermediate[4095+1719:0+1719] + a; end
12'd1720: begin if(a[1720]==1) 
	 		intermediate[4095+1720:0+1720] <= intermediate[4095+1720:0+1720] + a; end
12'd1721: begin if(a[1721]==1) 
	 		intermediate[4095+1721:0+1721] <= intermediate[4095+1721:0+1721] + a; end
12'd1722: begin if(a[1722]==1) 
	 		intermediate[4095+1722:0+1722] <= intermediate[4095+1722:0+1722] + a; end
12'd1723: begin if(a[1723]==1) 
	 		intermediate[4095+1723:0+1723] <= intermediate[4095+1723:0+1723] + a; end
12'd1724: begin if(a[1724]==1) 
	 		intermediate[4095+1724:0+1724] <= intermediate[4095+1724:0+1724] + a; end
12'd1725: begin if(a[1725]==1) 
	 		intermediate[4095+1725:0+1725] <= intermediate[4095+1725:0+1725] + a; end
12'd1726: begin if(a[1726]==1) 
	 		intermediate[4095+1726:0+1726] <= intermediate[4095+1726:0+1726] + a; end
12'd1727: begin if(a[1727]==1) 
	 		intermediate[4095+1727:0+1727] <= intermediate[4095+1727:0+1727] + a; end
12'd1728: begin if(a[1728]==1) 
	 		intermediate[4095+1728:0+1728] <= intermediate[4095+1728:0+1728] + a; end
12'd1729: begin if(a[1729]==1) 
	 		intermediate[4095+1729:0+1729] <= intermediate[4095+1729:0+1729] + a; end
12'd1730: begin if(a[1730]==1) 
	 		intermediate[4095+1730:0+1730] <= intermediate[4095+1730:0+1730] + a; end
12'd1731: begin if(a[1731]==1) 
	 		intermediate[4095+1731:0+1731] <= intermediate[4095+1731:0+1731] + a; end
12'd1732: begin if(a[1732]==1) 
	 		intermediate[4095+1732:0+1732] <= intermediate[4095+1732:0+1732] + a; end
12'd1733: begin if(a[1733]==1) 
	 		intermediate[4095+1733:0+1733] <= intermediate[4095+1733:0+1733] + a; end
12'd1734: begin if(a[1734]==1) 
	 		intermediate[4095+1734:0+1734] <= intermediate[4095+1734:0+1734] + a; end
12'd1735: begin if(a[1735]==1) 
	 		intermediate[4095+1735:0+1735] <= intermediate[4095+1735:0+1735] + a; end
12'd1736: begin if(a[1736]==1) 
	 		intermediate[4095+1736:0+1736] <= intermediate[4095+1736:0+1736] + a; end
12'd1737: begin if(a[1737]==1) 
	 		intermediate[4095+1737:0+1737] <= intermediate[4095+1737:0+1737] + a; end
12'd1738: begin if(a[1738]==1) 
	 		intermediate[4095+1738:0+1738] <= intermediate[4095+1738:0+1738] + a; end
12'd1739: begin if(a[1739]==1) 
	 		intermediate[4095+1739:0+1739] <= intermediate[4095+1739:0+1739] + a; end
12'd1740: begin if(a[1740]==1) 
	 		intermediate[4095+1740:0+1740] <= intermediate[4095+1740:0+1740] + a; end
12'd1741: begin if(a[1741]==1) 
	 		intermediate[4095+1741:0+1741] <= intermediate[4095+1741:0+1741] + a; end
12'd1742: begin if(a[1742]==1) 
	 		intermediate[4095+1742:0+1742] <= intermediate[4095+1742:0+1742] + a; end
12'd1743: begin if(a[1743]==1) 
	 		intermediate[4095+1743:0+1743] <= intermediate[4095+1743:0+1743] + a; end
12'd1744: begin if(a[1744]==1) 
	 		intermediate[4095+1744:0+1744] <= intermediate[4095+1744:0+1744] + a; end
12'd1745: begin if(a[1745]==1) 
	 		intermediate[4095+1745:0+1745] <= intermediate[4095+1745:0+1745] + a; end
12'd1746: begin if(a[1746]==1) 
	 		intermediate[4095+1746:0+1746] <= intermediate[4095+1746:0+1746] + a; end
12'd1747: begin if(a[1747]==1) 
	 		intermediate[4095+1747:0+1747] <= intermediate[4095+1747:0+1747] + a; end
12'd1748: begin if(a[1748]==1) 
	 		intermediate[4095+1748:0+1748] <= intermediate[4095+1748:0+1748] + a; end
12'd1749: begin if(a[1749]==1) 
	 		intermediate[4095+1749:0+1749] <= intermediate[4095+1749:0+1749] + a; end
12'd1750: begin if(a[1750]==1) 
	 		intermediate[4095+1750:0+1750] <= intermediate[4095+1750:0+1750] + a; end
12'd1751: begin if(a[1751]==1) 
	 		intermediate[4095+1751:0+1751] <= intermediate[4095+1751:0+1751] + a; end
12'd1752: begin if(a[1752]==1) 
	 		intermediate[4095+1752:0+1752] <= intermediate[4095+1752:0+1752] + a; end
12'd1753: begin if(a[1753]==1) 
	 		intermediate[4095+1753:0+1753] <= intermediate[4095+1753:0+1753] + a; end
12'd1754: begin if(a[1754]==1) 
	 		intermediate[4095+1754:0+1754] <= intermediate[4095+1754:0+1754] + a; end
12'd1755: begin if(a[1755]==1) 
	 		intermediate[4095+1755:0+1755] <= intermediate[4095+1755:0+1755] + a; end
12'd1756: begin if(a[1756]==1) 
	 		intermediate[4095+1756:0+1756] <= intermediate[4095+1756:0+1756] + a; end
12'd1757: begin if(a[1757]==1) 
	 		intermediate[4095+1757:0+1757] <= intermediate[4095+1757:0+1757] + a; end
12'd1758: begin if(a[1758]==1) 
	 		intermediate[4095+1758:0+1758] <= intermediate[4095+1758:0+1758] + a; end
12'd1759: begin if(a[1759]==1) 
	 		intermediate[4095+1759:0+1759] <= intermediate[4095+1759:0+1759] + a; end
12'd1760: begin if(a[1760]==1) 
	 		intermediate[4095+1760:0+1760] <= intermediate[4095+1760:0+1760] + a; end
12'd1761: begin if(a[1761]==1) 
	 		intermediate[4095+1761:0+1761] <= intermediate[4095+1761:0+1761] + a; end
12'd1762: begin if(a[1762]==1) 
	 		intermediate[4095+1762:0+1762] <= intermediate[4095+1762:0+1762] + a; end
12'd1763: begin if(a[1763]==1) 
	 		intermediate[4095+1763:0+1763] <= intermediate[4095+1763:0+1763] + a; end
12'd1764: begin if(a[1764]==1) 
	 		intermediate[4095+1764:0+1764] <= intermediate[4095+1764:0+1764] + a; end
12'd1765: begin if(a[1765]==1) 
	 		intermediate[4095+1765:0+1765] <= intermediate[4095+1765:0+1765] + a; end
12'd1766: begin if(a[1766]==1) 
	 		intermediate[4095+1766:0+1766] <= intermediate[4095+1766:0+1766] + a; end
12'd1767: begin if(a[1767]==1) 
	 		intermediate[4095+1767:0+1767] <= intermediate[4095+1767:0+1767] + a; end
12'd1768: begin if(a[1768]==1) 
	 		intermediate[4095+1768:0+1768] <= intermediate[4095+1768:0+1768] + a; end
12'd1769: begin if(a[1769]==1) 
	 		intermediate[4095+1769:0+1769] <= intermediate[4095+1769:0+1769] + a; end
12'd1770: begin if(a[1770]==1) 
	 		intermediate[4095+1770:0+1770] <= intermediate[4095+1770:0+1770] + a; end
12'd1771: begin if(a[1771]==1) 
	 		intermediate[4095+1771:0+1771] <= intermediate[4095+1771:0+1771] + a; end
12'd1772: begin if(a[1772]==1) 
	 		intermediate[4095+1772:0+1772] <= intermediate[4095+1772:0+1772] + a; end
12'd1773: begin if(a[1773]==1) 
	 		intermediate[4095+1773:0+1773] <= intermediate[4095+1773:0+1773] + a; end
12'd1774: begin if(a[1774]==1) 
	 		intermediate[4095+1774:0+1774] <= intermediate[4095+1774:0+1774] + a; end
12'd1775: begin if(a[1775]==1) 
	 		intermediate[4095+1775:0+1775] <= intermediate[4095+1775:0+1775] + a; end
12'd1776: begin if(a[1776]==1) 
	 		intermediate[4095+1776:0+1776] <= intermediate[4095+1776:0+1776] + a; end
12'd1777: begin if(a[1777]==1) 
	 		intermediate[4095+1777:0+1777] <= intermediate[4095+1777:0+1777] + a; end
12'd1778: begin if(a[1778]==1) 
	 		intermediate[4095+1778:0+1778] <= intermediate[4095+1778:0+1778] + a; end
12'd1779: begin if(a[1779]==1) 
	 		intermediate[4095+1779:0+1779] <= intermediate[4095+1779:0+1779] + a; end
12'd1780: begin if(a[1780]==1) 
	 		intermediate[4095+1780:0+1780] <= intermediate[4095+1780:0+1780] + a; end
12'd1781: begin if(a[1781]==1) 
	 		intermediate[4095+1781:0+1781] <= intermediate[4095+1781:0+1781] + a; end
12'd1782: begin if(a[1782]==1) 
	 		intermediate[4095+1782:0+1782] <= intermediate[4095+1782:0+1782] + a; end
12'd1783: begin if(a[1783]==1) 
	 		intermediate[4095+1783:0+1783] <= intermediate[4095+1783:0+1783] + a; end
12'd1784: begin if(a[1784]==1) 
	 		intermediate[4095+1784:0+1784] <= intermediate[4095+1784:0+1784] + a; end
12'd1785: begin if(a[1785]==1) 
	 		intermediate[4095+1785:0+1785] <= intermediate[4095+1785:0+1785] + a; end
12'd1786: begin if(a[1786]==1) 
	 		intermediate[4095+1786:0+1786] <= intermediate[4095+1786:0+1786] + a; end
12'd1787: begin if(a[1787]==1) 
	 		intermediate[4095+1787:0+1787] <= intermediate[4095+1787:0+1787] + a; end
12'd1788: begin if(a[1788]==1) 
	 		intermediate[4095+1788:0+1788] <= intermediate[4095+1788:0+1788] + a; end
12'd1789: begin if(a[1789]==1) 
	 		intermediate[4095+1789:0+1789] <= intermediate[4095+1789:0+1789] + a; end
12'd1790: begin if(a[1790]==1) 
	 		intermediate[4095+1790:0+1790] <= intermediate[4095+1790:0+1790] + a; end
12'd1791: begin if(a[1791]==1) 
	 		intermediate[4095+1791:0+1791] <= intermediate[4095+1791:0+1791] + a; end
12'd1792: begin if(a[1792]==1) 
	 		intermediate[4095+1792:0+1792] <= intermediate[4095+1792:0+1792] + a; end
12'd1793: begin if(a[1793]==1) 
	 		intermediate[4095+1793:0+1793] <= intermediate[4095+1793:0+1793] + a; end
12'd1794: begin if(a[1794]==1) 
	 		intermediate[4095+1794:0+1794] <= intermediate[4095+1794:0+1794] + a; end
12'd1795: begin if(a[1795]==1) 
	 		intermediate[4095+1795:0+1795] <= intermediate[4095+1795:0+1795] + a; end
12'd1796: begin if(a[1796]==1) 
	 		intermediate[4095+1796:0+1796] <= intermediate[4095+1796:0+1796] + a; end
12'd1797: begin if(a[1797]==1) 
	 		intermediate[4095+1797:0+1797] <= intermediate[4095+1797:0+1797] + a; end
12'd1798: begin if(a[1798]==1) 
	 		intermediate[4095+1798:0+1798] <= intermediate[4095+1798:0+1798] + a; end
12'd1799: begin if(a[1799]==1) 
	 		intermediate[4095+1799:0+1799] <= intermediate[4095+1799:0+1799] + a; end
12'd1800: begin if(a[1800]==1) 
	 		intermediate[4095+1800:0+1800] <= intermediate[4095+1800:0+1800] + a; end
12'd1801: begin if(a[1801]==1) 
	 		intermediate[4095+1801:0+1801] <= intermediate[4095+1801:0+1801] + a; end
12'd1802: begin if(a[1802]==1) 
	 		intermediate[4095+1802:0+1802] <= intermediate[4095+1802:0+1802] + a; end
12'd1803: begin if(a[1803]==1) 
	 		intermediate[4095+1803:0+1803] <= intermediate[4095+1803:0+1803] + a; end
12'd1804: begin if(a[1804]==1) 
	 		intermediate[4095+1804:0+1804] <= intermediate[4095+1804:0+1804] + a; end
12'd1805: begin if(a[1805]==1) 
	 		intermediate[4095+1805:0+1805] <= intermediate[4095+1805:0+1805] + a; end
12'd1806: begin if(a[1806]==1) 
	 		intermediate[4095+1806:0+1806] <= intermediate[4095+1806:0+1806] + a; end
12'd1807: begin if(a[1807]==1) 
	 		intermediate[4095+1807:0+1807] <= intermediate[4095+1807:0+1807] + a; end
12'd1808: begin if(a[1808]==1) 
	 		intermediate[4095+1808:0+1808] <= intermediate[4095+1808:0+1808] + a; end
12'd1809: begin if(a[1809]==1) 
	 		intermediate[4095+1809:0+1809] <= intermediate[4095+1809:0+1809] + a; end
12'd1810: begin if(a[1810]==1) 
	 		intermediate[4095+1810:0+1810] <= intermediate[4095+1810:0+1810] + a; end
12'd1811: begin if(a[1811]==1) 
	 		intermediate[4095+1811:0+1811] <= intermediate[4095+1811:0+1811] + a; end
12'd1812: begin if(a[1812]==1) 
	 		intermediate[4095+1812:0+1812] <= intermediate[4095+1812:0+1812] + a; end
12'd1813: begin if(a[1813]==1) 
	 		intermediate[4095+1813:0+1813] <= intermediate[4095+1813:0+1813] + a; end
12'd1814: begin if(a[1814]==1) 
	 		intermediate[4095+1814:0+1814] <= intermediate[4095+1814:0+1814] + a; end
12'd1815: begin if(a[1815]==1) 
	 		intermediate[4095+1815:0+1815] <= intermediate[4095+1815:0+1815] + a; end
12'd1816: begin if(a[1816]==1) 
	 		intermediate[4095+1816:0+1816] <= intermediate[4095+1816:0+1816] + a; end
12'd1817: begin if(a[1817]==1) 
	 		intermediate[4095+1817:0+1817] <= intermediate[4095+1817:0+1817] + a; end
12'd1818: begin if(a[1818]==1) 
	 		intermediate[4095+1818:0+1818] <= intermediate[4095+1818:0+1818] + a; end
12'd1819: begin if(a[1819]==1) 
	 		intermediate[4095+1819:0+1819] <= intermediate[4095+1819:0+1819] + a; end
12'd1820: begin if(a[1820]==1) 
	 		intermediate[4095+1820:0+1820] <= intermediate[4095+1820:0+1820] + a; end
12'd1821: begin if(a[1821]==1) 
	 		intermediate[4095+1821:0+1821] <= intermediate[4095+1821:0+1821] + a; end
12'd1822: begin if(a[1822]==1) 
	 		intermediate[4095+1822:0+1822] <= intermediate[4095+1822:0+1822] + a; end
12'd1823: begin if(a[1823]==1) 
	 		intermediate[4095+1823:0+1823] <= intermediate[4095+1823:0+1823] + a; end
12'd1824: begin if(a[1824]==1) 
	 		intermediate[4095+1824:0+1824] <= intermediate[4095+1824:0+1824] + a; end
12'd1825: begin if(a[1825]==1) 
	 		intermediate[4095+1825:0+1825] <= intermediate[4095+1825:0+1825] + a; end
12'd1826: begin if(a[1826]==1) 
	 		intermediate[4095+1826:0+1826] <= intermediate[4095+1826:0+1826] + a; end
12'd1827: begin if(a[1827]==1) 
	 		intermediate[4095+1827:0+1827] <= intermediate[4095+1827:0+1827] + a; end
12'd1828: begin if(a[1828]==1) 
	 		intermediate[4095+1828:0+1828] <= intermediate[4095+1828:0+1828] + a; end
12'd1829: begin if(a[1829]==1) 
	 		intermediate[4095+1829:0+1829] <= intermediate[4095+1829:0+1829] + a; end
12'd1830: begin if(a[1830]==1) 
	 		intermediate[4095+1830:0+1830] <= intermediate[4095+1830:0+1830] + a; end
12'd1831: begin if(a[1831]==1) 
	 		intermediate[4095+1831:0+1831] <= intermediate[4095+1831:0+1831] + a; end
12'd1832: begin if(a[1832]==1) 
	 		intermediate[4095+1832:0+1832] <= intermediate[4095+1832:0+1832] + a; end
12'd1833: begin if(a[1833]==1) 
	 		intermediate[4095+1833:0+1833] <= intermediate[4095+1833:0+1833] + a; end
12'd1834: begin if(a[1834]==1) 
	 		intermediate[4095+1834:0+1834] <= intermediate[4095+1834:0+1834] + a; end
12'd1835: begin if(a[1835]==1) 
	 		intermediate[4095+1835:0+1835] <= intermediate[4095+1835:0+1835] + a; end
12'd1836: begin if(a[1836]==1) 
	 		intermediate[4095+1836:0+1836] <= intermediate[4095+1836:0+1836] + a; end
12'd1837: begin if(a[1837]==1) 
	 		intermediate[4095+1837:0+1837] <= intermediate[4095+1837:0+1837] + a; end
12'd1838: begin if(a[1838]==1) 
	 		intermediate[4095+1838:0+1838] <= intermediate[4095+1838:0+1838] + a; end
12'd1839: begin if(a[1839]==1) 
	 		intermediate[4095+1839:0+1839] <= intermediate[4095+1839:0+1839] + a; end
12'd1840: begin if(a[1840]==1) 
	 		intermediate[4095+1840:0+1840] <= intermediate[4095+1840:0+1840] + a; end
12'd1841: begin if(a[1841]==1) 
	 		intermediate[4095+1841:0+1841] <= intermediate[4095+1841:0+1841] + a; end
12'd1842: begin if(a[1842]==1) 
	 		intermediate[4095+1842:0+1842] <= intermediate[4095+1842:0+1842] + a; end
12'd1843: begin if(a[1843]==1) 
	 		intermediate[4095+1843:0+1843] <= intermediate[4095+1843:0+1843] + a; end
12'd1844: begin if(a[1844]==1) 
	 		intermediate[4095+1844:0+1844] <= intermediate[4095+1844:0+1844] + a; end
12'd1845: begin if(a[1845]==1) 
	 		intermediate[4095+1845:0+1845] <= intermediate[4095+1845:0+1845] + a; end
12'd1846: begin if(a[1846]==1) 
	 		intermediate[4095+1846:0+1846] <= intermediate[4095+1846:0+1846] + a; end
12'd1847: begin if(a[1847]==1) 
	 		intermediate[4095+1847:0+1847] <= intermediate[4095+1847:0+1847] + a; end
12'd1848: begin if(a[1848]==1) 
	 		intermediate[4095+1848:0+1848] <= intermediate[4095+1848:0+1848] + a; end
12'd1849: begin if(a[1849]==1) 
	 		intermediate[4095+1849:0+1849] <= intermediate[4095+1849:0+1849] + a; end
12'd1850: begin if(a[1850]==1) 
	 		intermediate[4095+1850:0+1850] <= intermediate[4095+1850:0+1850] + a; end
12'd1851: begin if(a[1851]==1) 
	 		intermediate[4095+1851:0+1851] <= intermediate[4095+1851:0+1851] + a; end
12'd1852: begin if(a[1852]==1) 
	 		intermediate[4095+1852:0+1852] <= intermediate[4095+1852:0+1852] + a; end
12'd1853: begin if(a[1853]==1) 
	 		intermediate[4095+1853:0+1853] <= intermediate[4095+1853:0+1853] + a; end
12'd1854: begin if(a[1854]==1) 
	 		intermediate[4095+1854:0+1854] <= intermediate[4095+1854:0+1854] + a; end
12'd1855: begin if(a[1855]==1) 
	 		intermediate[4095+1855:0+1855] <= intermediate[4095+1855:0+1855] + a; end
12'd1856: begin if(a[1856]==1) 
	 		intermediate[4095+1856:0+1856] <= intermediate[4095+1856:0+1856] + a; end
12'd1857: begin if(a[1857]==1) 
	 		intermediate[4095+1857:0+1857] <= intermediate[4095+1857:0+1857] + a; end
12'd1858: begin if(a[1858]==1) 
	 		intermediate[4095+1858:0+1858] <= intermediate[4095+1858:0+1858] + a; end
12'd1859: begin if(a[1859]==1) 
	 		intermediate[4095+1859:0+1859] <= intermediate[4095+1859:0+1859] + a; end
12'd1860: begin if(a[1860]==1) 
	 		intermediate[4095+1860:0+1860] <= intermediate[4095+1860:0+1860] + a; end
12'd1861: begin if(a[1861]==1) 
	 		intermediate[4095+1861:0+1861] <= intermediate[4095+1861:0+1861] + a; end
12'd1862: begin if(a[1862]==1) 
	 		intermediate[4095+1862:0+1862] <= intermediate[4095+1862:0+1862] + a; end
12'd1863: begin if(a[1863]==1) 
	 		intermediate[4095+1863:0+1863] <= intermediate[4095+1863:0+1863] + a; end
12'd1864: begin if(a[1864]==1) 
	 		intermediate[4095+1864:0+1864] <= intermediate[4095+1864:0+1864] + a; end
12'd1865: begin if(a[1865]==1) 
	 		intermediate[4095+1865:0+1865] <= intermediate[4095+1865:0+1865] + a; end
12'd1866: begin if(a[1866]==1) 
	 		intermediate[4095+1866:0+1866] <= intermediate[4095+1866:0+1866] + a; end
12'd1867: begin if(a[1867]==1) 
	 		intermediate[4095+1867:0+1867] <= intermediate[4095+1867:0+1867] + a; end
12'd1868: begin if(a[1868]==1) 
	 		intermediate[4095+1868:0+1868] <= intermediate[4095+1868:0+1868] + a; end
12'd1869: begin if(a[1869]==1) 
	 		intermediate[4095+1869:0+1869] <= intermediate[4095+1869:0+1869] + a; end
12'd1870: begin if(a[1870]==1) 
	 		intermediate[4095+1870:0+1870] <= intermediate[4095+1870:0+1870] + a; end
12'd1871: begin if(a[1871]==1) 
	 		intermediate[4095+1871:0+1871] <= intermediate[4095+1871:0+1871] + a; end
12'd1872: begin if(a[1872]==1) 
	 		intermediate[4095+1872:0+1872] <= intermediate[4095+1872:0+1872] + a; end
12'd1873: begin if(a[1873]==1) 
	 		intermediate[4095+1873:0+1873] <= intermediate[4095+1873:0+1873] + a; end
12'd1874: begin if(a[1874]==1) 
	 		intermediate[4095+1874:0+1874] <= intermediate[4095+1874:0+1874] + a; end
12'd1875: begin if(a[1875]==1) 
	 		intermediate[4095+1875:0+1875] <= intermediate[4095+1875:0+1875] + a; end
12'd1876: begin if(a[1876]==1) 
	 		intermediate[4095+1876:0+1876] <= intermediate[4095+1876:0+1876] + a; end
12'd1877: begin if(a[1877]==1) 
	 		intermediate[4095+1877:0+1877] <= intermediate[4095+1877:0+1877] + a; end
12'd1878: begin if(a[1878]==1) 
	 		intermediate[4095+1878:0+1878] <= intermediate[4095+1878:0+1878] + a; end
12'd1879: begin if(a[1879]==1) 
	 		intermediate[4095+1879:0+1879] <= intermediate[4095+1879:0+1879] + a; end
12'd1880: begin if(a[1880]==1) 
	 		intermediate[4095+1880:0+1880] <= intermediate[4095+1880:0+1880] + a; end
12'd1881: begin if(a[1881]==1) 
	 		intermediate[4095+1881:0+1881] <= intermediate[4095+1881:0+1881] + a; end
12'd1882: begin if(a[1882]==1) 
	 		intermediate[4095+1882:0+1882] <= intermediate[4095+1882:0+1882] + a; end
12'd1883: begin if(a[1883]==1) 
	 		intermediate[4095+1883:0+1883] <= intermediate[4095+1883:0+1883] + a; end
12'd1884: begin if(a[1884]==1) 
	 		intermediate[4095+1884:0+1884] <= intermediate[4095+1884:0+1884] + a; end
12'd1885: begin if(a[1885]==1) 
	 		intermediate[4095+1885:0+1885] <= intermediate[4095+1885:0+1885] + a; end
12'd1886: begin if(a[1886]==1) 
	 		intermediate[4095+1886:0+1886] <= intermediate[4095+1886:0+1886] + a; end
12'd1887: begin if(a[1887]==1) 
	 		intermediate[4095+1887:0+1887] <= intermediate[4095+1887:0+1887] + a; end
12'd1888: begin if(a[1888]==1) 
	 		intermediate[4095+1888:0+1888] <= intermediate[4095+1888:0+1888] + a; end
12'd1889: begin if(a[1889]==1) 
	 		intermediate[4095+1889:0+1889] <= intermediate[4095+1889:0+1889] + a; end
12'd1890: begin if(a[1890]==1) 
	 		intermediate[4095+1890:0+1890] <= intermediate[4095+1890:0+1890] + a; end
12'd1891: begin if(a[1891]==1) 
	 		intermediate[4095+1891:0+1891] <= intermediate[4095+1891:0+1891] + a; end
12'd1892: begin if(a[1892]==1) 
	 		intermediate[4095+1892:0+1892] <= intermediate[4095+1892:0+1892] + a; end
12'd1893: begin if(a[1893]==1) 
	 		intermediate[4095+1893:0+1893] <= intermediate[4095+1893:0+1893] + a; end
12'd1894: begin if(a[1894]==1) 
	 		intermediate[4095+1894:0+1894] <= intermediate[4095+1894:0+1894] + a; end
12'd1895: begin if(a[1895]==1) 
	 		intermediate[4095+1895:0+1895] <= intermediate[4095+1895:0+1895] + a; end
12'd1896: begin if(a[1896]==1) 
	 		intermediate[4095+1896:0+1896] <= intermediate[4095+1896:0+1896] + a; end
12'd1897: begin if(a[1897]==1) 
	 		intermediate[4095+1897:0+1897] <= intermediate[4095+1897:0+1897] + a; end
12'd1898: begin if(a[1898]==1) 
	 		intermediate[4095+1898:0+1898] <= intermediate[4095+1898:0+1898] + a; end
12'd1899: begin if(a[1899]==1) 
	 		intermediate[4095+1899:0+1899] <= intermediate[4095+1899:0+1899] + a; end
12'd1900: begin if(a[1900]==1) 
	 		intermediate[4095+1900:0+1900] <= intermediate[4095+1900:0+1900] + a; end
12'd1901: begin if(a[1901]==1) 
	 		intermediate[4095+1901:0+1901] <= intermediate[4095+1901:0+1901] + a; end
12'd1902: begin if(a[1902]==1) 
	 		intermediate[4095+1902:0+1902] <= intermediate[4095+1902:0+1902] + a; end
12'd1903: begin if(a[1903]==1) 
	 		intermediate[4095+1903:0+1903] <= intermediate[4095+1903:0+1903] + a; end
12'd1904: begin if(a[1904]==1) 
	 		intermediate[4095+1904:0+1904] <= intermediate[4095+1904:0+1904] + a; end
12'd1905: begin if(a[1905]==1) 
	 		intermediate[4095+1905:0+1905] <= intermediate[4095+1905:0+1905] + a; end
12'd1906: begin if(a[1906]==1) 
	 		intermediate[4095+1906:0+1906] <= intermediate[4095+1906:0+1906] + a; end
12'd1907: begin if(a[1907]==1) 
	 		intermediate[4095+1907:0+1907] <= intermediate[4095+1907:0+1907] + a; end
12'd1908: begin if(a[1908]==1) 
	 		intermediate[4095+1908:0+1908] <= intermediate[4095+1908:0+1908] + a; end
12'd1909: begin if(a[1909]==1) 
	 		intermediate[4095+1909:0+1909] <= intermediate[4095+1909:0+1909] + a; end
12'd1910: begin if(a[1910]==1) 
	 		intermediate[4095+1910:0+1910] <= intermediate[4095+1910:0+1910] + a; end
12'd1911: begin if(a[1911]==1) 
	 		intermediate[4095+1911:0+1911] <= intermediate[4095+1911:0+1911] + a; end
12'd1912: begin if(a[1912]==1) 
	 		intermediate[4095+1912:0+1912] <= intermediate[4095+1912:0+1912] + a; end
12'd1913: begin if(a[1913]==1) 
	 		intermediate[4095+1913:0+1913] <= intermediate[4095+1913:0+1913] + a; end
12'd1914: begin if(a[1914]==1) 
	 		intermediate[4095+1914:0+1914] <= intermediate[4095+1914:0+1914] + a; end
12'd1915: begin if(a[1915]==1) 
	 		intermediate[4095+1915:0+1915] <= intermediate[4095+1915:0+1915] + a; end
12'd1916: begin if(a[1916]==1) 
	 		intermediate[4095+1916:0+1916] <= intermediate[4095+1916:0+1916] + a; end
12'd1917: begin if(a[1917]==1) 
	 		intermediate[4095+1917:0+1917] <= intermediate[4095+1917:0+1917] + a; end
12'd1918: begin if(a[1918]==1) 
	 		intermediate[4095+1918:0+1918] <= intermediate[4095+1918:0+1918] + a; end
12'd1919: begin if(a[1919]==1) 
	 		intermediate[4095+1919:0+1919] <= intermediate[4095+1919:0+1919] + a; end
12'd1920: begin if(a[1920]==1) 
	 		intermediate[4095+1920:0+1920] <= intermediate[4095+1920:0+1920] + a; end
12'd1921: begin if(a[1921]==1) 
	 		intermediate[4095+1921:0+1921] <= intermediate[4095+1921:0+1921] + a; end
12'd1922: begin if(a[1922]==1) 
	 		intermediate[4095+1922:0+1922] <= intermediate[4095+1922:0+1922] + a; end
12'd1923: begin if(a[1923]==1) 
	 		intermediate[4095+1923:0+1923] <= intermediate[4095+1923:0+1923] + a; end
12'd1924: begin if(a[1924]==1) 
	 		intermediate[4095+1924:0+1924] <= intermediate[4095+1924:0+1924] + a; end
12'd1925: begin if(a[1925]==1) 
	 		intermediate[4095+1925:0+1925] <= intermediate[4095+1925:0+1925] + a; end
12'd1926: begin if(a[1926]==1) 
	 		intermediate[4095+1926:0+1926] <= intermediate[4095+1926:0+1926] + a; end
12'd1927: begin if(a[1927]==1) 
	 		intermediate[4095+1927:0+1927] <= intermediate[4095+1927:0+1927] + a; end
12'd1928: begin if(a[1928]==1) 
	 		intermediate[4095+1928:0+1928] <= intermediate[4095+1928:0+1928] + a; end
12'd1929: begin if(a[1929]==1) 
	 		intermediate[4095+1929:0+1929] <= intermediate[4095+1929:0+1929] + a; end
12'd1930: begin if(a[1930]==1) 
	 		intermediate[4095+1930:0+1930] <= intermediate[4095+1930:0+1930] + a; end
12'd1931: begin if(a[1931]==1) 
	 		intermediate[4095+1931:0+1931] <= intermediate[4095+1931:0+1931] + a; end
12'd1932: begin if(a[1932]==1) 
	 		intermediate[4095+1932:0+1932] <= intermediate[4095+1932:0+1932] + a; end
12'd1933: begin if(a[1933]==1) 
	 		intermediate[4095+1933:0+1933] <= intermediate[4095+1933:0+1933] + a; end
12'd1934: begin if(a[1934]==1) 
	 		intermediate[4095+1934:0+1934] <= intermediate[4095+1934:0+1934] + a; end
12'd1935: begin if(a[1935]==1) 
	 		intermediate[4095+1935:0+1935] <= intermediate[4095+1935:0+1935] + a; end
12'd1936: begin if(a[1936]==1) 
	 		intermediate[4095+1936:0+1936] <= intermediate[4095+1936:0+1936] + a; end
12'd1937: begin if(a[1937]==1) 
	 		intermediate[4095+1937:0+1937] <= intermediate[4095+1937:0+1937] + a; end
12'd1938: begin if(a[1938]==1) 
	 		intermediate[4095+1938:0+1938] <= intermediate[4095+1938:0+1938] + a; end
12'd1939: begin if(a[1939]==1) 
	 		intermediate[4095+1939:0+1939] <= intermediate[4095+1939:0+1939] + a; end
12'd1940: begin if(a[1940]==1) 
	 		intermediate[4095+1940:0+1940] <= intermediate[4095+1940:0+1940] + a; end
12'd1941: begin if(a[1941]==1) 
	 		intermediate[4095+1941:0+1941] <= intermediate[4095+1941:0+1941] + a; end
12'd1942: begin if(a[1942]==1) 
	 		intermediate[4095+1942:0+1942] <= intermediate[4095+1942:0+1942] + a; end
12'd1943: begin if(a[1943]==1) 
	 		intermediate[4095+1943:0+1943] <= intermediate[4095+1943:0+1943] + a; end
12'd1944: begin if(a[1944]==1) 
	 		intermediate[4095+1944:0+1944] <= intermediate[4095+1944:0+1944] + a; end
12'd1945: begin if(a[1945]==1) 
	 		intermediate[4095+1945:0+1945] <= intermediate[4095+1945:0+1945] + a; end
12'd1946: begin if(a[1946]==1) 
	 		intermediate[4095+1946:0+1946] <= intermediate[4095+1946:0+1946] + a; end
12'd1947: begin if(a[1947]==1) 
	 		intermediate[4095+1947:0+1947] <= intermediate[4095+1947:0+1947] + a; end
12'd1948: begin if(a[1948]==1) 
	 		intermediate[4095+1948:0+1948] <= intermediate[4095+1948:0+1948] + a; end
12'd1949: begin if(a[1949]==1) 
	 		intermediate[4095+1949:0+1949] <= intermediate[4095+1949:0+1949] + a; end
12'd1950: begin if(a[1950]==1) 
	 		intermediate[4095+1950:0+1950] <= intermediate[4095+1950:0+1950] + a; end
12'd1951: begin if(a[1951]==1) 
	 		intermediate[4095+1951:0+1951] <= intermediate[4095+1951:0+1951] + a; end
12'd1952: begin if(a[1952]==1) 
	 		intermediate[4095+1952:0+1952] <= intermediate[4095+1952:0+1952] + a; end
12'd1953: begin if(a[1953]==1) 
	 		intermediate[4095+1953:0+1953] <= intermediate[4095+1953:0+1953] + a; end
12'd1954: begin if(a[1954]==1) 
	 		intermediate[4095+1954:0+1954] <= intermediate[4095+1954:0+1954] + a; end
12'd1955: begin if(a[1955]==1) 
	 		intermediate[4095+1955:0+1955] <= intermediate[4095+1955:0+1955] + a; end
12'd1956: begin if(a[1956]==1) 
	 		intermediate[4095+1956:0+1956] <= intermediate[4095+1956:0+1956] + a; end
12'd1957: begin if(a[1957]==1) 
	 		intermediate[4095+1957:0+1957] <= intermediate[4095+1957:0+1957] + a; end
12'd1958: begin if(a[1958]==1) 
	 		intermediate[4095+1958:0+1958] <= intermediate[4095+1958:0+1958] + a; end
12'd1959: begin if(a[1959]==1) 
	 		intermediate[4095+1959:0+1959] <= intermediate[4095+1959:0+1959] + a; end
12'd1960: begin if(a[1960]==1) 
	 		intermediate[4095+1960:0+1960] <= intermediate[4095+1960:0+1960] + a; end
12'd1961: begin if(a[1961]==1) 
	 		intermediate[4095+1961:0+1961] <= intermediate[4095+1961:0+1961] + a; end
12'd1962: begin if(a[1962]==1) 
	 		intermediate[4095+1962:0+1962] <= intermediate[4095+1962:0+1962] + a; end
12'd1963: begin if(a[1963]==1) 
	 		intermediate[4095+1963:0+1963] <= intermediate[4095+1963:0+1963] + a; end
12'd1964: begin if(a[1964]==1) 
	 		intermediate[4095+1964:0+1964] <= intermediate[4095+1964:0+1964] + a; end
12'd1965: begin if(a[1965]==1) 
	 		intermediate[4095+1965:0+1965] <= intermediate[4095+1965:0+1965] + a; end
12'd1966: begin if(a[1966]==1) 
	 		intermediate[4095+1966:0+1966] <= intermediate[4095+1966:0+1966] + a; end
12'd1967: begin if(a[1967]==1) 
	 		intermediate[4095+1967:0+1967] <= intermediate[4095+1967:0+1967] + a; end
12'd1968: begin if(a[1968]==1) 
	 		intermediate[4095+1968:0+1968] <= intermediate[4095+1968:0+1968] + a; end
12'd1969: begin if(a[1969]==1) 
	 		intermediate[4095+1969:0+1969] <= intermediate[4095+1969:0+1969] + a; end
12'd1970: begin if(a[1970]==1) 
	 		intermediate[4095+1970:0+1970] <= intermediate[4095+1970:0+1970] + a; end
12'd1971: begin if(a[1971]==1) 
	 		intermediate[4095+1971:0+1971] <= intermediate[4095+1971:0+1971] + a; end
12'd1972: begin if(a[1972]==1) 
	 		intermediate[4095+1972:0+1972] <= intermediate[4095+1972:0+1972] + a; end
12'd1973: begin if(a[1973]==1) 
	 		intermediate[4095+1973:0+1973] <= intermediate[4095+1973:0+1973] + a; end
12'd1974: begin if(a[1974]==1) 
	 		intermediate[4095+1974:0+1974] <= intermediate[4095+1974:0+1974] + a; end
12'd1975: begin if(a[1975]==1) 
	 		intermediate[4095+1975:0+1975] <= intermediate[4095+1975:0+1975] + a; end
12'd1976: begin if(a[1976]==1) 
	 		intermediate[4095+1976:0+1976] <= intermediate[4095+1976:0+1976] + a; end
12'd1977: begin if(a[1977]==1) 
	 		intermediate[4095+1977:0+1977] <= intermediate[4095+1977:0+1977] + a; end
12'd1978: begin if(a[1978]==1) 
	 		intermediate[4095+1978:0+1978] <= intermediate[4095+1978:0+1978] + a; end
12'd1979: begin if(a[1979]==1) 
	 		intermediate[4095+1979:0+1979] <= intermediate[4095+1979:0+1979] + a; end
12'd1980: begin if(a[1980]==1) 
	 		intermediate[4095+1980:0+1980] <= intermediate[4095+1980:0+1980] + a; end
12'd1981: begin if(a[1981]==1) 
	 		intermediate[4095+1981:0+1981] <= intermediate[4095+1981:0+1981] + a; end
12'd1982: begin if(a[1982]==1) 
	 		intermediate[4095+1982:0+1982] <= intermediate[4095+1982:0+1982] + a; end
12'd1983: begin if(a[1983]==1) 
	 		intermediate[4095+1983:0+1983] <= intermediate[4095+1983:0+1983] + a; end
12'd1984: begin if(a[1984]==1) 
	 		intermediate[4095+1984:0+1984] <= intermediate[4095+1984:0+1984] + a; end
12'd1985: begin if(a[1985]==1) 
	 		intermediate[4095+1985:0+1985] <= intermediate[4095+1985:0+1985] + a; end
12'd1986: begin if(a[1986]==1) 
	 		intermediate[4095+1986:0+1986] <= intermediate[4095+1986:0+1986] + a; end
12'd1987: begin if(a[1987]==1) 
	 		intermediate[4095+1987:0+1987] <= intermediate[4095+1987:0+1987] + a; end
12'd1988: begin if(a[1988]==1) 
	 		intermediate[4095+1988:0+1988] <= intermediate[4095+1988:0+1988] + a; end
12'd1989: begin if(a[1989]==1) 
	 		intermediate[4095+1989:0+1989] <= intermediate[4095+1989:0+1989] + a; end
12'd1990: begin if(a[1990]==1) 
	 		intermediate[4095+1990:0+1990] <= intermediate[4095+1990:0+1990] + a; end
12'd1991: begin if(a[1991]==1) 
	 		intermediate[4095+1991:0+1991] <= intermediate[4095+1991:0+1991] + a; end
12'd1992: begin if(a[1992]==1) 
	 		intermediate[4095+1992:0+1992] <= intermediate[4095+1992:0+1992] + a; end
12'd1993: begin if(a[1993]==1) 
	 		intermediate[4095+1993:0+1993] <= intermediate[4095+1993:0+1993] + a; end
12'd1994: begin if(a[1994]==1) 
	 		intermediate[4095+1994:0+1994] <= intermediate[4095+1994:0+1994] + a; end
12'd1995: begin if(a[1995]==1) 
	 		intermediate[4095+1995:0+1995] <= intermediate[4095+1995:0+1995] + a; end
12'd1996: begin if(a[1996]==1) 
	 		intermediate[4095+1996:0+1996] <= intermediate[4095+1996:0+1996] + a; end
12'd1997: begin if(a[1997]==1) 
	 		intermediate[4095+1997:0+1997] <= intermediate[4095+1997:0+1997] + a; end
12'd1998: begin if(a[1998]==1) 
	 		intermediate[4095+1998:0+1998] <= intermediate[4095+1998:0+1998] + a; end
12'd1999: begin if(a[1999]==1) 
	 		intermediate[4095+1999:0+1999] <= intermediate[4095+1999:0+1999] + a; end
12'd2000: begin if(a[2000]==1) 
	 		intermediate[4095+2000:0+2000] <= intermediate[4095+2000:0+2000] + a; end
12'd2001: begin if(a[2001]==1) 
	 		intermediate[4095+2001:0+2001] <= intermediate[4095+2001:0+2001] + a; end
12'd2002: begin if(a[2002]==1) 
	 		intermediate[4095+2002:0+2002] <= intermediate[4095+2002:0+2002] + a; end
12'd2003: begin if(a[2003]==1) 
	 		intermediate[4095+2003:0+2003] <= intermediate[4095+2003:0+2003] + a; end
12'd2004: begin if(a[2004]==1) 
	 		intermediate[4095+2004:0+2004] <= intermediate[4095+2004:0+2004] + a; end
12'd2005: begin if(a[2005]==1) 
	 		intermediate[4095+2005:0+2005] <= intermediate[4095+2005:0+2005] + a; end
12'd2006: begin if(a[2006]==1) 
	 		intermediate[4095+2006:0+2006] <= intermediate[4095+2006:0+2006] + a; end
12'd2007: begin if(a[2007]==1) 
	 		intermediate[4095+2007:0+2007] <= intermediate[4095+2007:0+2007] + a; end
12'd2008: begin if(a[2008]==1) 
	 		intermediate[4095+2008:0+2008] <= intermediate[4095+2008:0+2008] + a; end
12'd2009: begin if(a[2009]==1) 
	 		intermediate[4095+2009:0+2009] <= intermediate[4095+2009:0+2009] + a; end
12'd2010: begin if(a[2010]==1) 
	 		intermediate[4095+2010:0+2010] <= intermediate[4095+2010:0+2010] + a; end
12'd2011: begin if(a[2011]==1) 
	 		intermediate[4095+2011:0+2011] <= intermediate[4095+2011:0+2011] + a; end
12'd2012: begin if(a[2012]==1) 
	 		intermediate[4095+2012:0+2012] <= intermediate[4095+2012:0+2012] + a; end
12'd2013: begin if(a[2013]==1) 
	 		intermediate[4095+2013:0+2013] <= intermediate[4095+2013:0+2013] + a; end
12'd2014: begin if(a[2014]==1) 
	 		intermediate[4095+2014:0+2014] <= intermediate[4095+2014:0+2014] + a; end
12'd2015: begin if(a[2015]==1) 
	 		intermediate[4095+2015:0+2015] <= intermediate[4095+2015:0+2015] + a; end
12'd2016: begin if(a[2016]==1) 
	 		intermediate[4095+2016:0+2016] <= intermediate[4095+2016:0+2016] + a; end
12'd2017: begin if(a[2017]==1) 
	 		intermediate[4095+2017:0+2017] <= intermediate[4095+2017:0+2017] + a; end
12'd2018: begin if(a[2018]==1) 
	 		intermediate[4095+2018:0+2018] <= intermediate[4095+2018:0+2018] + a; end
12'd2019: begin if(a[2019]==1) 
	 		intermediate[4095+2019:0+2019] <= intermediate[4095+2019:0+2019] + a; end
12'd2020: begin if(a[2020]==1) 
	 		intermediate[4095+2020:0+2020] <= intermediate[4095+2020:0+2020] + a; end
12'd2021: begin if(a[2021]==1) 
	 		intermediate[4095+2021:0+2021] <= intermediate[4095+2021:0+2021] + a; end
12'd2022: begin if(a[2022]==1) 
	 		intermediate[4095+2022:0+2022] <= intermediate[4095+2022:0+2022] + a; end
12'd2023: begin if(a[2023]==1) 
	 		intermediate[4095+2023:0+2023] <= intermediate[4095+2023:0+2023] + a; end
12'd2024: begin if(a[2024]==1) 
	 		intermediate[4095+2024:0+2024] <= intermediate[4095+2024:0+2024] + a; end
12'd2025: begin if(a[2025]==1) 
	 		intermediate[4095+2025:0+2025] <= intermediate[4095+2025:0+2025] + a; end
12'd2026: begin if(a[2026]==1) 
	 		intermediate[4095+2026:0+2026] <= intermediate[4095+2026:0+2026] + a; end
12'd2027: begin if(a[2027]==1) 
	 		intermediate[4095+2027:0+2027] <= intermediate[4095+2027:0+2027] + a; end
12'd2028: begin if(a[2028]==1) 
	 		intermediate[4095+2028:0+2028] <= intermediate[4095+2028:0+2028] + a; end
12'd2029: begin if(a[2029]==1) 
	 		intermediate[4095+2029:0+2029] <= intermediate[4095+2029:0+2029] + a; end
12'd2030: begin if(a[2030]==1) 
	 		intermediate[4095+2030:0+2030] <= intermediate[4095+2030:0+2030] + a; end
12'd2031: begin if(a[2031]==1) 
	 		intermediate[4095+2031:0+2031] <= intermediate[4095+2031:0+2031] + a; end
12'd2032: begin if(a[2032]==1) 
	 		intermediate[4095+2032:0+2032] <= intermediate[4095+2032:0+2032] + a; end
12'd2033: begin if(a[2033]==1) 
	 		intermediate[4095+2033:0+2033] <= intermediate[4095+2033:0+2033] + a; end
12'd2034: begin if(a[2034]==1) 
	 		intermediate[4095+2034:0+2034] <= intermediate[4095+2034:0+2034] + a; end
12'd2035: begin if(a[2035]==1) 
	 		intermediate[4095+2035:0+2035] <= intermediate[4095+2035:0+2035] + a; end
12'd2036: begin if(a[2036]==1) 
	 		intermediate[4095+2036:0+2036] <= intermediate[4095+2036:0+2036] + a; end
12'd2037: begin if(a[2037]==1) 
	 		intermediate[4095+2037:0+2037] <= intermediate[4095+2037:0+2037] + a; end
12'd2038: begin if(a[2038]==1) 
	 		intermediate[4095+2038:0+2038] <= intermediate[4095+2038:0+2038] + a; end
12'd2039: begin if(a[2039]==1) 
	 		intermediate[4095+2039:0+2039] <= intermediate[4095+2039:0+2039] + a; end
12'd2040: begin if(a[2040]==1) 
	 		intermediate[4095+2040:0+2040] <= intermediate[4095+2040:0+2040] + a; end
12'd2041: begin if(a[2041]==1) 
	 		intermediate[4095+2041:0+2041] <= intermediate[4095+2041:0+2041] + a; end
12'd2042: begin if(a[2042]==1) 
	 		intermediate[4095+2042:0+2042] <= intermediate[4095+2042:0+2042] + a; end
12'd2043: begin if(a[2043]==1) 
	 		intermediate[4095+2043:0+2043] <= intermediate[4095+2043:0+2043] + a; end
12'd2044: begin if(a[2044]==1) 
	 		intermediate[4095+2044:0+2044] <= intermediate[4095+2044:0+2044] + a; end
12'd2045: begin if(a[2045]==1) 
	 		intermediate[4095+2045:0+2045] <= intermediate[4095+2045:0+2045] + a; end
12'd2046: begin if(a[2046]==1) 
	 		intermediate[4095+2046:0+2046] <= intermediate[4095+2046:0+2046] + a; end
12'd2047: begin if(a[2047]==1) 
	 		intermediate[4095+2047:0+2047] <= intermediate[4095+2047:0+2047] + a; end
12'd2048: begin if(a[2048]==1) 
	 		intermediate[4095+2048:0+2048] <= intermediate[4095+2048:0+2048] + a; end
12'd2049: begin if(a[2049]==1) 
	 		intermediate[4095+2049:0+2049] <= intermediate[4095+2049:0+2049] + a; end
12'd2050: begin if(a[2050]==1) 
	 		intermediate[4095+2050:0+2050] <= intermediate[4095+2050:0+2050] + a; end
12'd2051: begin if(a[2051]==1) 
	 		intermediate[4095+2051:0+2051] <= intermediate[4095+2051:0+2051] + a; end
12'd2052: begin if(a[2052]==1) 
	 		intermediate[4095+2052:0+2052] <= intermediate[4095+2052:0+2052] + a; end
12'd2053: begin if(a[2053]==1) 
	 		intermediate[4095+2053:0+2053] <= intermediate[4095+2053:0+2053] + a; end
12'd2054: begin if(a[2054]==1) 
	 		intermediate[4095+2054:0+2054] <= intermediate[4095+2054:0+2054] + a; end
12'd2055: begin if(a[2055]==1) 
	 		intermediate[4095+2055:0+2055] <= intermediate[4095+2055:0+2055] + a; end
12'd2056: begin if(a[2056]==1) 
	 		intermediate[4095+2056:0+2056] <= intermediate[4095+2056:0+2056] + a; end
12'd2057: begin if(a[2057]==1) 
	 		intermediate[4095+2057:0+2057] <= intermediate[4095+2057:0+2057] + a; end
12'd2058: begin if(a[2058]==1) 
	 		intermediate[4095+2058:0+2058] <= intermediate[4095+2058:0+2058] + a; end
12'd2059: begin if(a[2059]==1) 
	 		intermediate[4095+2059:0+2059] <= intermediate[4095+2059:0+2059] + a; end
12'd2060: begin if(a[2060]==1) 
	 		intermediate[4095+2060:0+2060] <= intermediate[4095+2060:0+2060] + a; end
12'd2061: begin if(a[2061]==1) 
	 		intermediate[4095+2061:0+2061] <= intermediate[4095+2061:0+2061] + a; end
12'd2062: begin if(a[2062]==1) 
	 		intermediate[4095+2062:0+2062] <= intermediate[4095+2062:0+2062] + a; end
12'd2063: begin if(a[2063]==1) 
	 		intermediate[4095+2063:0+2063] <= intermediate[4095+2063:0+2063] + a; end
12'd2064: begin if(a[2064]==1) 
	 		intermediate[4095+2064:0+2064] <= intermediate[4095+2064:0+2064] + a; end
12'd2065: begin if(a[2065]==1) 
	 		intermediate[4095+2065:0+2065] <= intermediate[4095+2065:0+2065] + a; end
12'd2066: begin if(a[2066]==1) 
	 		intermediate[4095+2066:0+2066] <= intermediate[4095+2066:0+2066] + a; end
12'd2067: begin if(a[2067]==1) 
	 		intermediate[4095+2067:0+2067] <= intermediate[4095+2067:0+2067] + a; end
12'd2068: begin if(a[2068]==1) 
	 		intermediate[4095+2068:0+2068] <= intermediate[4095+2068:0+2068] + a; end
12'd2069: begin if(a[2069]==1) 
	 		intermediate[4095+2069:0+2069] <= intermediate[4095+2069:0+2069] + a; end
12'd2070: begin if(a[2070]==1) 
	 		intermediate[4095+2070:0+2070] <= intermediate[4095+2070:0+2070] + a; end
12'd2071: begin if(a[2071]==1) 
	 		intermediate[4095+2071:0+2071] <= intermediate[4095+2071:0+2071] + a; end
12'd2072: begin if(a[2072]==1) 
	 		intermediate[4095+2072:0+2072] <= intermediate[4095+2072:0+2072] + a; end
12'd2073: begin if(a[2073]==1) 
	 		intermediate[4095+2073:0+2073] <= intermediate[4095+2073:0+2073] + a; end
12'd2074: begin if(a[2074]==1) 
	 		intermediate[4095+2074:0+2074] <= intermediate[4095+2074:0+2074] + a; end
12'd2075: begin if(a[2075]==1) 
	 		intermediate[4095+2075:0+2075] <= intermediate[4095+2075:0+2075] + a; end
12'd2076: begin if(a[2076]==1) 
	 		intermediate[4095+2076:0+2076] <= intermediate[4095+2076:0+2076] + a; end
12'd2077: begin if(a[2077]==1) 
	 		intermediate[4095+2077:0+2077] <= intermediate[4095+2077:0+2077] + a; end
12'd2078: begin if(a[2078]==1) 
	 		intermediate[4095+2078:0+2078] <= intermediate[4095+2078:0+2078] + a; end
12'd2079: begin if(a[2079]==1) 
	 		intermediate[4095+2079:0+2079] <= intermediate[4095+2079:0+2079] + a; end
12'd2080: begin if(a[2080]==1) 
	 		intermediate[4095+2080:0+2080] <= intermediate[4095+2080:0+2080] + a; end
12'd2081: begin if(a[2081]==1) 
	 		intermediate[4095+2081:0+2081] <= intermediate[4095+2081:0+2081] + a; end
12'd2082: begin if(a[2082]==1) 
	 		intermediate[4095+2082:0+2082] <= intermediate[4095+2082:0+2082] + a; end
12'd2083: begin if(a[2083]==1) 
	 		intermediate[4095+2083:0+2083] <= intermediate[4095+2083:0+2083] + a; end
12'd2084: begin if(a[2084]==1) 
	 		intermediate[4095+2084:0+2084] <= intermediate[4095+2084:0+2084] + a; end
12'd2085: begin if(a[2085]==1) 
	 		intermediate[4095+2085:0+2085] <= intermediate[4095+2085:0+2085] + a; end
12'd2086: begin if(a[2086]==1) 
	 		intermediate[4095+2086:0+2086] <= intermediate[4095+2086:0+2086] + a; end
12'd2087: begin if(a[2087]==1) 
	 		intermediate[4095+2087:0+2087] <= intermediate[4095+2087:0+2087] + a; end
12'd2088: begin if(a[2088]==1) 
	 		intermediate[4095+2088:0+2088] <= intermediate[4095+2088:0+2088] + a; end
12'd2089: begin if(a[2089]==1) 
	 		intermediate[4095+2089:0+2089] <= intermediate[4095+2089:0+2089] + a; end
12'd2090: begin if(a[2090]==1) 
	 		intermediate[4095+2090:0+2090] <= intermediate[4095+2090:0+2090] + a; end
12'd2091: begin if(a[2091]==1) 
	 		intermediate[4095+2091:0+2091] <= intermediate[4095+2091:0+2091] + a; end
12'd2092: begin if(a[2092]==1) 
	 		intermediate[4095+2092:0+2092] <= intermediate[4095+2092:0+2092] + a; end
12'd2093: begin if(a[2093]==1) 
	 		intermediate[4095+2093:0+2093] <= intermediate[4095+2093:0+2093] + a; end
12'd2094: begin if(a[2094]==1) 
	 		intermediate[4095+2094:0+2094] <= intermediate[4095+2094:0+2094] + a; end
12'd2095: begin if(a[2095]==1) 
	 		intermediate[4095+2095:0+2095] <= intermediate[4095+2095:0+2095] + a; end
12'd2096: begin if(a[2096]==1) 
	 		intermediate[4095+2096:0+2096] <= intermediate[4095+2096:0+2096] + a; end
12'd2097: begin if(a[2097]==1) 
	 		intermediate[4095+2097:0+2097] <= intermediate[4095+2097:0+2097] + a; end
12'd2098: begin if(a[2098]==1) 
	 		intermediate[4095+2098:0+2098] <= intermediate[4095+2098:0+2098] + a; end
12'd2099: begin if(a[2099]==1) 
	 		intermediate[4095+2099:0+2099] <= intermediate[4095+2099:0+2099] + a; end
12'd2100: begin if(a[2100]==1) 
	 		intermediate[4095+2100:0+2100] <= intermediate[4095+2100:0+2100] + a; end
12'd2101: begin if(a[2101]==1) 
	 		intermediate[4095+2101:0+2101] <= intermediate[4095+2101:0+2101] + a; end
12'd2102: begin if(a[2102]==1) 
	 		intermediate[4095+2102:0+2102] <= intermediate[4095+2102:0+2102] + a; end
12'd2103: begin if(a[2103]==1) 
	 		intermediate[4095+2103:0+2103] <= intermediate[4095+2103:0+2103] + a; end
12'd2104: begin if(a[2104]==1) 
	 		intermediate[4095+2104:0+2104] <= intermediate[4095+2104:0+2104] + a; end
12'd2105: begin if(a[2105]==1) 
	 		intermediate[4095+2105:0+2105] <= intermediate[4095+2105:0+2105] + a; end
12'd2106: begin if(a[2106]==1) 
	 		intermediate[4095+2106:0+2106] <= intermediate[4095+2106:0+2106] + a; end
12'd2107: begin if(a[2107]==1) 
	 		intermediate[4095+2107:0+2107] <= intermediate[4095+2107:0+2107] + a; end
12'd2108: begin if(a[2108]==1) 
	 		intermediate[4095+2108:0+2108] <= intermediate[4095+2108:0+2108] + a; end
12'd2109: begin if(a[2109]==1) 
	 		intermediate[4095+2109:0+2109] <= intermediate[4095+2109:0+2109] + a; end
12'd2110: begin if(a[2110]==1) 
	 		intermediate[4095+2110:0+2110] <= intermediate[4095+2110:0+2110] + a; end
12'd2111: begin if(a[2111]==1) 
	 		intermediate[4095+2111:0+2111] <= intermediate[4095+2111:0+2111] + a; end
12'd2112: begin if(a[2112]==1) 
	 		intermediate[4095+2112:0+2112] <= intermediate[4095+2112:0+2112] + a; end
12'd2113: begin if(a[2113]==1) 
	 		intermediate[4095+2113:0+2113] <= intermediate[4095+2113:0+2113] + a; end
12'd2114: begin if(a[2114]==1) 
	 		intermediate[4095+2114:0+2114] <= intermediate[4095+2114:0+2114] + a; end
12'd2115: begin if(a[2115]==1) 
	 		intermediate[4095+2115:0+2115] <= intermediate[4095+2115:0+2115] + a; end
12'd2116: begin if(a[2116]==1) 
	 		intermediate[4095+2116:0+2116] <= intermediate[4095+2116:0+2116] + a; end
12'd2117: begin if(a[2117]==1) 
	 		intermediate[4095+2117:0+2117] <= intermediate[4095+2117:0+2117] + a; end
12'd2118: begin if(a[2118]==1) 
	 		intermediate[4095+2118:0+2118] <= intermediate[4095+2118:0+2118] + a; end
12'd2119: begin if(a[2119]==1) 
	 		intermediate[4095+2119:0+2119] <= intermediate[4095+2119:0+2119] + a; end
12'd2120: begin if(a[2120]==1) 
	 		intermediate[4095+2120:0+2120] <= intermediate[4095+2120:0+2120] + a; end
12'd2121: begin if(a[2121]==1) 
	 		intermediate[4095+2121:0+2121] <= intermediate[4095+2121:0+2121] + a; end
12'd2122: begin if(a[2122]==1) 
	 		intermediate[4095+2122:0+2122] <= intermediate[4095+2122:0+2122] + a; end
12'd2123: begin if(a[2123]==1) 
	 		intermediate[4095+2123:0+2123] <= intermediate[4095+2123:0+2123] + a; end
12'd2124: begin if(a[2124]==1) 
	 		intermediate[4095+2124:0+2124] <= intermediate[4095+2124:0+2124] + a; end
12'd2125: begin if(a[2125]==1) 
	 		intermediate[4095+2125:0+2125] <= intermediate[4095+2125:0+2125] + a; end
12'd2126: begin if(a[2126]==1) 
	 		intermediate[4095+2126:0+2126] <= intermediate[4095+2126:0+2126] + a; end
12'd2127: begin if(a[2127]==1) 
	 		intermediate[4095+2127:0+2127] <= intermediate[4095+2127:0+2127] + a; end
12'd2128: begin if(a[2128]==1) 
	 		intermediate[4095+2128:0+2128] <= intermediate[4095+2128:0+2128] + a; end
12'd2129: begin if(a[2129]==1) 
	 		intermediate[4095+2129:0+2129] <= intermediate[4095+2129:0+2129] + a; end
12'd2130: begin if(a[2130]==1) 
	 		intermediate[4095+2130:0+2130] <= intermediate[4095+2130:0+2130] + a; end
12'd2131: begin if(a[2131]==1) 
	 		intermediate[4095+2131:0+2131] <= intermediate[4095+2131:0+2131] + a; end
12'd2132: begin if(a[2132]==1) 
	 		intermediate[4095+2132:0+2132] <= intermediate[4095+2132:0+2132] + a; end
12'd2133: begin if(a[2133]==1) 
	 		intermediate[4095+2133:0+2133] <= intermediate[4095+2133:0+2133] + a; end
12'd2134: begin if(a[2134]==1) 
	 		intermediate[4095+2134:0+2134] <= intermediate[4095+2134:0+2134] + a; end
12'd2135: begin if(a[2135]==1) 
	 		intermediate[4095+2135:0+2135] <= intermediate[4095+2135:0+2135] + a; end
12'd2136: begin if(a[2136]==1) 
	 		intermediate[4095+2136:0+2136] <= intermediate[4095+2136:0+2136] + a; end
12'd2137: begin if(a[2137]==1) 
	 		intermediate[4095+2137:0+2137] <= intermediate[4095+2137:0+2137] + a; end
12'd2138: begin if(a[2138]==1) 
	 		intermediate[4095+2138:0+2138] <= intermediate[4095+2138:0+2138] + a; end
12'd2139: begin if(a[2139]==1) 
	 		intermediate[4095+2139:0+2139] <= intermediate[4095+2139:0+2139] + a; end
12'd2140: begin if(a[2140]==1) 
	 		intermediate[4095+2140:0+2140] <= intermediate[4095+2140:0+2140] + a; end
12'd2141: begin if(a[2141]==1) 
	 		intermediate[4095+2141:0+2141] <= intermediate[4095+2141:0+2141] + a; end
12'd2142: begin if(a[2142]==1) 
	 		intermediate[4095+2142:0+2142] <= intermediate[4095+2142:0+2142] + a; end
12'd2143: begin if(a[2143]==1) 
	 		intermediate[4095+2143:0+2143] <= intermediate[4095+2143:0+2143] + a; end
12'd2144: begin if(a[2144]==1) 
	 		intermediate[4095+2144:0+2144] <= intermediate[4095+2144:0+2144] + a; end
12'd2145: begin if(a[2145]==1) 
	 		intermediate[4095+2145:0+2145] <= intermediate[4095+2145:0+2145] + a; end
12'd2146: begin if(a[2146]==1) 
	 		intermediate[4095+2146:0+2146] <= intermediate[4095+2146:0+2146] + a; end
12'd2147: begin if(a[2147]==1) 
	 		intermediate[4095+2147:0+2147] <= intermediate[4095+2147:0+2147] + a; end
12'd2148: begin if(a[2148]==1) 
	 		intermediate[4095+2148:0+2148] <= intermediate[4095+2148:0+2148] + a; end
12'd2149: begin if(a[2149]==1) 
	 		intermediate[4095+2149:0+2149] <= intermediate[4095+2149:0+2149] + a; end
12'd2150: begin if(a[2150]==1) 
	 		intermediate[4095+2150:0+2150] <= intermediate[4095+2150:0+2150] + a; end
12'd2151: begin if(a[2151]==1) 
	 		intermediate[4095+2151:0+2151] <= intermediate[4095+2151:0+2151] + a; end
12'd2152: begin if(a[2152]==1) 
	 		intermediate[4095+2152:0+2152] <= intermediate[4095+2152:0+2152] + a; end
12'd2153: begin if(a[2153]==1) 
	 		intermediate[4095+2153:0+2153] <= intermediate[4095+2153:0+2153] + a; end
12'd2154: begin if(a[2154]==1) 
	 		intermediate[4095+2154:0+2154] <= intermediate[4095+2154:0+2154] + a; end
12'd2155: begin if(a[2155]==1) 
	 		intermediate[4095+2155:0+2155] <= intermediate[4095+2155:0+2155] + a; end
12'd2156: begin if(a[2156]==1) 
	 		intermediate[4095+2156:0+2156] <= intermediate[4095+2156:0+2156] + a; end
12'd2157: begin if(a[2157]==1) 
	 		intermediate[4095+2157:0+2157] <= intermediate[4095+2157:0+2157] + a; end
12'd2158: begin if(a[2158]==1) 
	 		intermediate[4095+2158:0+2158] <= intermediate[4095+2158:0+2158] + a; end
12'd2159: begin if(a[2159]==1) 
	 		intermediate[4095+2159:0+2159] <= intermediate[4095+2159:0+2159] + a; end
12'd2160: begin if(a[2160]==1) 
	 		intermediate[4095+2160:0+2160] <= intermediate[4095+2160:0+2160] + a; end
12'd2161: begin if(a[2161]==1) 
	 		intermediate[4095+2161:0+2161] <= intermediate[4095+2161:0+2161] + a; end
12'd2162: begin if(a[2162]==1) 
	 		intermediate[4095+2162:0+2162] <= intermediate[4095+2162:0+2162] + a; end
12'd2163: begin if(a[2163]==1) 
	 		intermediate[4095+2163:0+2163] <= intermediate[4095+2163:0+2163] + a; end
12'd2164: begin if(a[2164]==1) 
	 		intermediate[4095+2164:0+2164] <= intermediate[4095+2164:0+2164] + a; end
12'd2165: begin if(a[2165]==1) 
	 		intermediate[4095+2165:0+2165] <= intermediate[4095+2165:0+2165] + a; end
12'd2166: begin if(a[2166]==1) 
	 		intermediate[4095+2166:0+2166] <= intermediate[4095+2166:0+2166] + a; end
12'd2167: begin if(a[2167]==1) 
	 		intermediate[4095+2167:0+2167] <= intermediate[4095+2167:0+2167] + a; end
12'd2168: begin if(a[2168]==1) 
	 		intermediate[4095+2168:0+2168] <= intermediate[4095+2168:0+2168] + a; end
12'd2169: begin if(a[2169]==1) 
	 		intermediate[4095+2169:0+2169] <= intermediate[4095+2169:0+2169] + a; end
12'd2170: begin if(a[2170]==1) 
	 		intermediate[4095+2170:0+2170] <= intermediate[4095+2170:0+2170] + a; end
12'd2171: begin if(a[2171]==1) 
	 		intermediate[4095+2171:0+2171] <= intermediate[4095+2171:0+2171] + a; end
12'd2172: begin if(a[2172]==1) 
	 		intermediate[4095+2172:0+2172] <= intermediate[4095+2172:0+2172] + a; end
12'd2173: begin if(a[2173]==1) 
	 		intermediate[4095+2173:0+2173] <= intermediate[4095+2173:0+2173] + a; end
12'd2174: begin if(a[2174]==1) 
	 		intermediate[4095+2174:0+2174] <= intermediate[4095+2174:0+2174] + a; end
12'd2175: begin if(a[2175]==1) 
	 		intermediate[4095+2175:0+2175] <= intermediate[4095+2175:0+2175] + a; end
12'd2176: begin if(a[2176]==1) 
	 		intermediate[4095+2176:0+2176] <= intermediate[4095+2176:0+2176] + a; end
12'd2177: begin if(a[2177]==1) 
	 		intermediate[4095+2177:0+2177] <= intermediate[4095+2177:0+2177] + a; end
12'd2178: begin if(a[2178]==1) 
	 		intermediate[4095+2178:0+2178] <= intermediate[4095+2178:0+2178] + a; end
12'd2179: begin if(a[2179]==1) 
	 		intermediate[4095+2179:0+2179] <= intermediate[4095+2179:0+2179] + a; end
12'd2180: begin if(a[2180]==1) 
	 		intermediate[4095+2180:0+2180] <= intermediate[4095+2180:0+2180] + a; end
12'd2181: begin if(a[2181]==1) 
	 		intermediate[4095+2181:0+2181] <= intermediate[4095+2181:0+2181] + a; end
12'd2182: begin if(a[2182]==1) 
	 		intermediate[4095+2182:0+2182] <= intermediate[4095+2182:0+2182] + a; end
12'd2183: begin if(a[2183]==1) 
	 		intermediate[4095+2183:0+2183] <= intermediate[4095+2183:0+2183] + a; end
12'd2184: begin if(a[2184]==1) 
	 		intermediate[4095+2184:0+2184] <= intermediate[4095+2184:0+2184] + a; end
12'd2185: begin if(a[2185]==1) 
	 		intermediate[4095+2185:0+2185] <= intermediate[4095+2185:0+2185] + a; end
12'd2186: begin if(a[2186]==1) 
	 		intermediate[4095+2186:0+2186] <= intermediate[4095+2186:0+2186] + a; end
12'd2187: begin if(a[2187]==1) 
	 		intermediate[4095+2187:0+2187] <= intermediate[4095+2187:0+2187] + a; end
12'd2188: begin if(a[2188]==1) 
	 		intermediate[4095+2188:0+2188] <= intermediate[4095+2188:0+2188] + a; end
12'd2189: begin if(a[2189]==1) 
	 		intermediate[4095+2189:0+2189] <= intermediate[4095+2189:0+2189] + a; end
12'd2190: begin if(a[2190]==1) 
	 		intermediate[4095+2190:0+2190] <= intermediate[4095+2190:0+2190] + a; end
12'd2191: begin if(a[2191]==1) 
	 		intermediate[4095+2191:0+2191] <= intermediate[4095+2191:0+2191] + a; end
12'd2192: begin if(a[2192]==1) 
	 		intermediate[4095+2192:0+2192] <= intermediate[4095+2192:0+2192] + a; end
12'd2193: begin if(a[2193]==1) 
	 		intermediate[4095+2193:0+2193] <= intermediate[4095+2193:0+2193] + a; end
12'd2194: begin if(a[2194]==1) 
	 		intermediate[4095+2194:0+2194] <= intermediate[4095+2194:0+2194] + a; end
12'd2195: begin if(a[2195]==1) 
	 		intermediate[4095+2195:0+2195] <= intermediate[4095+2195:0+2195] + a; end
12'd2196: begin if(a[2196]==1) 
	 		intermediate[4095+2196:0+2196] <= intermediate[4095+2196:0+2196] + a; end
12'd2197: begin if(a[2197]==1) 
	 		intermediate[4095+2197:0+2197] <= intermediate[4095+2197:0+2197] + a; end
12'd2198: begin if(a[2198]==1) 
	 		intermediate[4095+2198:0+2198] <= intermediate[4095+2198:0+2198] + a; end
12'd2199: begin if(a[2199]==1) 
	 		intermediate[4095+2199:0+2199] <= intermediate[4095+2199:0+2199] + a; end
12'd2200: begin if(a[2200]==1) 
	 		intermediate[4095+2200:0+2200] <= intermediate[4095+2200:0+2200] + a; end
12'd2201: begin if(a[2201]==1) 
	 		intermediate[4095+2201:0+2201] <= intermediate[4095+2201:0+2201] + a; end
12'd2202: begin if(a[2202]==1) 
	 		intermediate[4095+2202:0+2202] <= intermediate[4095+2202:0+2202] + a; end
12'd2203: begin if(a[2203]==1) 
	 		intermediate[4095+2203:0+2203] <= intermediate[4095+2203:0+2203] + a; end
12'd2204: begin if(a[2204]==1) 
	 		intermediate[4095+2204:0+2204] <= intermediate[4095+2204:0+2204] + a; end
12'd2205: begin if(a[2205]==1) 
	 		intermediate[4095+2205:0+2205] <= intermediate[4095+2205:0+2205] + a; end
12'd2206: begin if(a[2206]==1) 
	 		intermediate[4095+2206:0+2206] <= intermediate[4095+2206:0+2206] + a; end
12'd2207: begin if(a[2207]==1) 
	 		intermediate[4095+2207:0+2207] <= intermediate[4095+2207:0+2207] + a; end
12'd2208: begin if(a[2208]==1) 
	 		intermediate[4095+2208:0+2208] <= intermediate[4095+2208:0+2208] + a; end
12'd2209: begin if(a[2209]==1) 
	 		intermediate[4095+2209:0+2209] <= intermediate[4095+2209:0+2209] + a; end
12'd2210: begin if(a[2210]==1) 
	 		intermediate[4095+2210:0+2210] <= intermediate[4095+2210:0+2210] + a; end
12'd2211: begin if(a[2211]==1) 
	 		intermediate[4095+2211:0+2211] <= intermediate[4095+2211:0+2211] + a; end
12'd2212: begin if(a[2212]==1) 
	 		intermediate[4095+2212:0+2212] <= intermediate[4095+2212:0+2212] + a; end
12'd2213: begin if(a[2213]==1) 
	 		intermediate[4095+2213:0+2213] <= intermediate[4095+2213:0+2213] + a; end
12'd2214: begin if(a[2214]==1) 
	 		intermediate[4095+2214:0+2214] <= intermediate[4095+2214:0+2214] + a; end
12'd2215: begin if(a[2215]==1) 
	 		intermediate[4095+2215:0+2215] <= intermediate[4095+2215:0+2215] + a; end
12'd2216: begin if(a[2216]==1) 
	 		intermediate[4095+2216:0+2216] <= intermediate[4095+2216:0+2216] + a; end
12'd2217: begin if(a[2217]==1) 
	 		intermediate[4095+2217:0+2217] <= intermediate[4095+2217:0+2217] + a; end
12'd2218: begin if(a[2218]==1) 
	 		intermediate[4095+2218:0+2218] <= intermediate[4095+2218:0+2218] + a; end
12'd2219: begin if(a[2219]==1) 
	 		intermediate[4095+2219:0+2219] <= intermediate[4095+2219:0+2219] + a; end
12'd2220: begin if(a[2220]==1) 
	 		intermediate[4095+2220:0+2220] <= intermediate[4095+2220:0+2220] + a; end
12'd2221: begin if(a[2221]==1) 
	 		intermediate[4095+2221:0+2221] <= intermediate[4095+2221:0+2221] + a; end
12'd2222: begin if(a[2222]==1) 
	 		intermediate[4095+2222:0+2222] <= intermediate[4095+2222:0+2222] + a; end
12'd2223: begin if(a[2223]==1) 
	 		intermediate[4095+2223:0+2223] <= intermediate[4095+2223:0+2223] + a; end
12'd2224: begin if(a[2224]==1) 
	 		intermediate[4095+2224:0+2224] <= intermediate[4095+2224:0+2224] + a; end
12'd2225: begin if(a[2225]==1) 
	 		intermediate[4095+2225:0+2225] <= intermediate[4095+2225:0+2225] + a; end
12'd2226: begin if(a[2226]==1) 
	 		intermediate[4095+2226:0+2226] <= intermediate[4095+2226:0+2226] + a; end
12'd2227: begin if(a[2227]==1) 
	 		intermediate[4095+2227:0+2227] <= intermediate[4095+2227:0+2227] + a; end
12'd2228: begin if(a[2228]==1) 
	 		intermediate[4095+2228:0+2228] <= intermediate[4095+2228:0+2228] + a; end
12'd2229: begin if(a[2229]==1) 
	 		intermediate[4095+2229:0+2229] <= intermediate[4095+2229:0+2229] + a; end
12'd2230: begin if(a[2230]==1) 
	 		intermediate[4095+2230:0+2230] <= intermediate[4095+2230:0+2230] + a; end
12'd2231: begin if(a[2231]==1) 
	 		intermediate[4095+2231:0+2231] <= intermediate[4095+2231:0+2231] + a; end
12'd2232: begin if(a[2232]==1) 
	 		intermediate[4095+2232:0+2232] <= intermediate[4095+2232:0+2232] + a; end
12'd2233: begin if(a[2233]==1) 
	 		intermediate[4095+2233:0+2233] <= intermediate[4095+2233:0+2233] + a; end
12'd2234: begin if(a[2234]==1) 
	 		intermediate[4095+2234:0+2234] <= intermediate[4095+2234:0+2234] + a; end
12'd2235: begin if(a[2235]==1) 
	 		intermediate[4095+2235:0+2235] <= intermediate[4095+2235:0+2235] + a; end
12'd2236: begin if(a[2236]==1) 
	 		intermediate[4095+2236:0+2236] <= intermediate[4095+2236:0+2236] + a; end
12'd2237: begin if(a[2237]==1) 
	 		intermediate[4095+2237:0+2237] <= intermediate[4095+2237:0+2237] + a; end
12'd2238: begin if(a[2238]==1) 
	 		intermediate[4095+2238:0+2238] <= intermediate[4095+2238:0+2238] + a; end
12'd2239: begin if(a[2239]==1) 
	 		intermediate[4095+2239:0+2239] <= intermediate[4095+2239:0+2239] + a; end
12'd2240: begin if(a[2240]==1) 
	 		intermediate[4095+2240:0+2240] <= intermediate[4095+2240:0+2240] + a; end
12'd2241: begin if(a[2241]==1) 
	 		intermediate[4095+2241:0+2241] <= intermediate[4095+2241:0+2241] + a; end
12'd2242: begin if(a[2242]==1) 
	 		intermediate[4095+2242:0+2242] <= intermediate[4095+2242:0+2242] + a; end
12'd2243: begin if(a[2243]==1) 
	 		intermediate[4095+2243:0+2243] <= intermediate[4095+2243:0+2243] + a; end
12'd2244: begin if(a[2244]==1) 
	 		intermediate[4095+2244:0+2244] <= intermediate[4095+2244:0+2244] + a; end
12'd2245: begin if(a[2245]==1) 
	 		intermediate[4095+2245:0+2245] <= intermediate[4095+2245:0+2245] + a; end
12'd2246: begin if(a[2246]==1) 
	 		intermediate[4095+2246:0+2246] <= intermediate[4095+2246:0+2246] + a; end
12'd2247: begin if(a[2247]==1) 
	 		intermediate[4095+2247:0+2247] <= intermediate[4095+2247:0+2247] + a; end
12'd2248: begin if(a[2248]==1) 
	 		intermediate[4095+2248:0+2248] <= intermediate[4095+2248:0+2248] + a; end
12'd2249: begin if(a[2249]==1) 
	 		intermediate[4095+2249:0+2249] <= intermediate[4095+2249:0+2249] + a; end
12'd2250: begin if(a[2250]==1) 
	 		intermediate[4095+2250:0+2250] <= intermediate[4095+2250:0+2250] + a; end
12'd2251: begin if(a[2251]==1) 
	 		intermediate[4095+2251:0+2251] <= intermediate[4095+2251:0+2251] + a; end
12'd2252: begin if(a[2252]==1) 
	 		intermediate[4095+2252:0+2252] <= intermediate[4095+2252:0+2252] + a; end
12'd2253: begin if(a[2253]==1) 
	 		intermediate[4095+2253:0+2253] <= intermediate[4095+2253:0+2253] + a; end
12'd2254: begin if(a[2254]==1) 
	 		intermediate[4095+2254:0+2254] <= intermediate[4095+2254:0+2254] + a; end
12'd2255: begin if(a[2255]==1) 
	 		intermediate[4095+2255:0+2255] <= intermediate[4095+2255:0+2255] + a; end
12'd2256: begin if(a[2256]==1) 
	 		intermediate[4095+2256:0+2256] <= intermediate[4095+2256:0+2256] + a; end
12'd2257: begin if(a[2257]==1) 
	 		intermediate[4095+2257:0+2257] <= intermediate[4095+2257:0+2257] + a; end
12'd2258: begin if(a[2258]==1) 
	 		intermediate[4095+2258:0+2258] <= intermediate[4095+2258:0+2258] + a; end
12'd2259: begin if(a[2259]==1) 
	 		intermediate[4095+2259:0+2259] <= intermediate[4095+2259:0+2259] + a; end
12'd2260: begin if(a[2260]==1) 
	 		intermediate[4095+2260:0+2260] <= intermediate[4095+2260:0+2260] + a; end
12'd2261: begin if(a[2261]==1) 
	 		intermediate[4095+2261:0+2261] <= intermediate[4095+2261:0+2261] + a; end
12'd2262: begin if(a[2262]==1) 
	 		intermediate[4095+2262:0+2262] <= intermediate[4095+2262:0+2262] + a; end
12'd2263: begin if(a[2263]==1) 
	 		intermediate[4095+2263:0+2263] <= intermediate[4095+2263:0+2263] + a; end
12'd2264: begin if(a[2264]==1) 
	 		intermediate[4095+2264:0+2264] <= intermediate[4095+2264:0+2264] + a; end
12'd2265: begin if(a[2265]==1) 
	 		intermediate[4095+2265:0+2265] <= intermediate[4095+2265:0+2265] + a; end
12'd2266: begin if(a[2266]==1) 
	 		intermediate[4095+2266:0+2266] <= intermediate[4095+2266:0+2266] + a; end
12'd2267: begin if(a[2267]==1) 
	 		intermediate[4095+2267:0+2267] <= intermediate[4095+2267:0+2267] + a; end
12'd2268: begin if(a[2268]==1) 
	 		intermediate[4095+2268:0+2268] <= intermediate[4095+2268:0+2268] + a; end
12'd2269: begin if(a[2269]==1) 
	 		intermediate[4095+2269:0+2269] <= intermediate[4095+2269:0+2269] + a; end
12'd2270: begin if(a[2270]==1) 
	 		intermediate[4095+2270:0+2270] <= intermediate[4095+2270:0+2270] + a; end
12'd2271: begin if(a[2271]==1) 
	 		intermediate[4095+2271:0+2271] <= intermediate[4095+2271:0+2271] + a; end
12'd2272: begin if(a[2272]==1) 
	 		intermediate[4095+2272:0+2272] <= intermediate[4095+2272:0+2272] + a; end
12'd2273: begin if(a[2273]==1) 
	 		intermediate[4095+2273:0+2273] <= intermediate[4095+2273:0+2273] + a; end
12'd2274: begin if(a[2274]==1) 
	 		intermediate[4095+2274:0+2274] <= intermediate[4095+2274:0+2274] + a; end
12'd2275: begin if(a[2275]==1) 
	 		intermediate[4095+2275:0+2275] <= intermediate[4095+2275:0+2275] + a; end
12'd2276: begin if(a[2276]==1) 
	 		intermediate[4095+2276:0+2276] <= intermediate[4095+2276:0+2276] + a; end
12'd2277: begin if(a[2277]==1) 
	 		intermediate[4095+2277:0+2277] <= intermediate[4095+2277:0+2277] + a; end
12'd2278: begin if(a[2278]==1) 
	 		intermediate[4095+2278:0+2278] <= intermediate[4095+2278:0+2278] + a; end
12'd2279: begin if(a[2279]==1) 
	 		intermediate[4095+2279:0+2279] <= intermediate[4095+2279:0+2279] + a; end
12'd2280: begin if(a[2280]==1) 
	 		intermediate[4095+2280:0+2280] <= intermediate[4095+2280:0+2280] + a; end
12'd2281: begin if(a[2281]==1) 
	 		intermediate[4095+2281:0+2281] <= intermediate[4095+2281:0+2281] + a; end
12'd2282: begin if(a[2282]==1) 
	 		intermediate[4095+2282:0+2282] <= intermediate[4095+2282:0+2282] + a; end
12'd2283: begin if(a[2283]==1) 
	 		intermediate[4095+2283:0+2283] <= intermediate[4095+2283:0+2283] + a; end
12'd2284: begin if(a[2284]==1) 
	 		intermediate[4095+2284:0+2284] <= intermediate[4095+2284:0+2284] + a; end
12'd2285: begin if(a[2285]==1) 
	 		intermediate[4095+2285:0+2285] <= intermediate[4095+2285:0+2285] + a; end
12'd2286: begin if(a[2286]==1) 
	 		intermediate[4095+2286:0+2286] <= intermediate[4095+2286:0+2286] + a; end
12'd2287: begin if(a[2287]==1) 
	 		intermediate[4095+2287:0+2287] <= intermediate[4095+2287:0+2287] + a; end
12'd2288: begin if(a[2288]==1) 
	 		intermediate[4095+2288:0+2288] <= intermediate[4095+2288:0+2288] + a; end
12'd2289: begin if(a[2289]==1) 
	 		intermediate[4095+2289:0+2289] <= intermediate[4095+2289:0+2289] + a; end
12'd2290: begin if(a[2290]==1) 
	 		intermediate[4095+2290:0+2290] <= intermediate[4095+2290:0+2290] + a; end
12'd2291: begin if(a[2291]==1) 
	 		intermediate[4095+2291:0+2291] <= intermediate[4095+2291:0+2291] + a; end
12'd2292: begin if(a[2292]==1) 
	 		intermediate[4095+2292:0+2292] <= intermediate[4095+2292:0+2292] + a; end
12'd2293: begin if(a[2293]==1) 
	 		intermediate[4095+2293:0+2293] <= intermediate[4095+2293:0+2293] + a; end
12'd2294: begin if(a[2294]==1) 
	 		intermediate[4095+2294:0+2294] <= intermediate[4095+2294:0+2294] + a; end
12'd2295: begin if(a[2295]==1) 
	 		intermediate[4095+2295:0+2295] <= intermediate[4095+2295:0+2295] + a; end
12'd2296: begin if(a[2296]==1) 
	 		intermediate[4095+2296:0+2296] <= intermediate[4095+2296:0+2296] + a; end
12'd2297: begin if(a[2297]==1) 
	 		intermediate[4095+2297:0+2297] <= intermediate[4095+2297:0+2297] + a; end
12'd2298: begin if(a[2298]==1) 
	 		intermediate[4095+2298:0+2298] <= intermediate[4095+2298:0+2298] + a; end
12'd2299: begin if(a[2299]==1) 
	 		intermediate[4095+2299:0+2299] <= intermediate[4095+2299:0+2299] + a; end
12'd2300: begin if(a[2300]==1) 
	 		intermediate[4095+2300:0+2300] <= intermediate[4095+2300:0+2300] + a; end
12'd2301: begin if(a[2301]==1) 
	 		intermediate[4095+2301:0+2301] <= intermediate[4095+2301:0+2301] + a; end
12'd2302: begin if(a[2302]==1) 
	 		intermediate[4095+2302:0+2302] <= intermediate[4095+2302:0+2302] + a; end
12'd2303: begin if(a[2303]==1) 
	 		intermediate[4095+2303:0+2303] <= intermediate[4095+2303:0+2303] + a; end
12'd2304: begin if(a[2304]==1) 
	 		intermediate[4095+2304:0+2304] <= intermediate[4095+2304:0+2304] + a; end
12'd2305: begin if(a[2305]==1) 
	 		intermediate[4095+2305:0+2305] <= intermediate[4095+2305:0+2305] + a; end
12'd2306: begin if(a[2306]==1) 
	 		intermediate[4095+2306:0+2306] <= intermediate[4095+2306:0+2306] + a; end
12'd2307: begin if(a[2307]==1) 
	 		intermediate[4095+2307:0+2307] <= intermediate[4095+2307:0+2307] + a; end
12'd2308: begin if(a[2308]==1) 
	 		intermediate[4095+2308:0+2308] <= intermediate[4095+2308:0+2308] + a; end
12'd2309: begin if(a[2309]==1) 
	 		intermediate[4095+2309:0+2309] <= intermediate[4095+2309:0+2309] + a; end
12'd2310: begin if(a[2310]==1) 
	 		intermediate[4095+2310:0+2310] <= intermediate[4095+2310:0+2310] + a; end
12'd2311: begin if(a[2311]==1) 
	 		intermediate[4095+2311:0+2311] <= intermediate[4095+2311:0+2311] + a; end
12'd2312: begin if(a[2312]==1) 
	 		intermediate[4095+2312:0+2312] <= intermediate[4095+2312:0+2312] + a; end
12'd2313: begin if(a[2313]==1) 
	 		intermediate[4095+2313:0+2313] <= intermediate[4095+2313:0+2313] + a; end
12'd2314: begin if(a[2314]==1) 
	 		intermediate[4095+2314:0+2314] <= intermediate[4095+2314:0+2314] + a; end
12'd2315: begin if(a[2315]==1) 
	 		intermediate[4095+2315:0+2315] <= intermediate[4095+2315:0+2315] + a; end
12'd2316: begin if(a[2316]==1) 
	 		intermediate[4095+2316:0+2316] <= intermediate[4095+2316:0+2316] + a; end
12'd2317: begin if(a[2317]==1) 
	 		intermediate[4095+2317:0+2317] <= intermediate[4095+2317:0+2317] + a; end
12'd2318: begin if(a[2318]==1) 
	 		intermediate[4095+2318:0+2318] <= intermediate[4095+2318:0+2318] + a; end
12'd2319: begin if(a[2319]==1) 
	 		intermediate[4095+2319:0+2319] <= intermediate[4095+2319:0+2319] + a; end
12'd2320: begin if(a[2320]==1) 
	 		intermediate[4095+2320:0+2320] <= intermediate[4095+2320:0+2320] + a; end
12'd2321: begin if(a[2321]==1) 
	 		intermediate[4095+2321:0+2321] <= intermediate[4095+2321:0+2321] + a; end
12'd2322: begin if(a[2322]==1) 
	 		intermediate[4095+2322:0+2322] <= intermediate[4095+2322:0+2322] + a; end
12'd2323: begin if(a[2323]==1) 
	 		intermediate[4095+2323:0+2323] <= intermediate[4095+2323:0+2323] + a; end
12'd2324: begin if(a[2324]==1) 
	 		intermediate[4095+2324:0+2324] <= intermediate[4095+2324:0+2324] + a; end
12'd2325: begin if(a[2325]==1) 
	 		intermediate[4095+2325:0+2325] <= intermediate[4095+2325:0+2325] + a; end
12'd2326: begin if(a[2326]==1) 
	 		intermediate[4095+2326:0+2326] <= intermediate[4095+2326:0+2326] + a; end
12'd2327: begin if(a[2327]==1) 
	 		intermediate[4095+2327:0+2327] <= intermediate[4095+2327:0+2327] + a; end
12'd2328: begin if(a[2328]==1) 
	 		intermediate[4095+2328:0+2328] <= intermediate[4095+2328:0+2328] + a; end
12'd2329: begin if(a[2329]==1) 
	 		intermediate[4095+2329:0+2329] <= intermediate[4095+2329:0+2329] + a; end
12'd2330: begin if(a[2330]==1) 
	 		intermediate[4095+2330:0+2330] <= intermediate[4095+2330:0+2330] + a; end
12'd2331: begin if(a[2331]==1) 
	 		intermediate[4095+2331:0+2331] <= intermediate[4095+2331:0+2331] + a; end
12'd2332: begin if(a[2332]==1) 
	 		intermediate[4095+2332:0+2332] <= intermediate[4095+2332:0+2332] + a; end
12'd2333: begin if(a[2333]==1) 
	 		intermediate[4095+2333:0+2333] <= intermediate[4095+2333:0+2333] + a; end
12'd2334: begin if(a[2334]==1) 
	 		intermediate[4095+2334:0+2334] <= intermediate[4095+2334:0+2334] + a; end
12'd2335: begin if(a[2335]==1) 
	 		intermediate[4095+2335:0+2335] <= intermediate[4095+2335:0+2335] + a; end
12'd2336: begin if(a[2336]==1) 
	 		intermediate[4095+2336:0+2336] <= intermediate[4095+2336:0+2336] + a; end
12'd2337: begin if(a[2337]==1) 
	 		intermediate[4095+2337:0+2337] <= intermediate[4095+2337:0+2337] + a; end
12'd2338: begin if(a[2338]==1) 
	 		intermediate[4095+2338:0+2338] <= intermediate[4095+2338:0+2338] + a; end
12'd2339: begin if(a[2339]==1) 
	 		intermediate[4095+2339:0+2339] <= intermediate[4095+2339:0+2339] + a; end
12'd2340: begin if(a[2340]==1) 
	 		intermediate[4095+2340:0+2340] <= intermediate[4095+2340:0+2340] + a; end
12'd2341: begin if(a[2341]==1) 
	 		intermediate[4095+2341:0+2341] <= intermediate[4095+2341:0+2341] + a; end
12'd2342: begin if(a[2342]==1) 
	 		intermediate[4095+2342:0+2342] <= intermediate[4095+2342:0+2342] + a; end
12'd2343: begin if(a[2343]==1) 
	 		intermediate[4095+2343:0+2343] <= intermediate[4095+2343:0+2343] + a; end
12'd2344: begin if(a[2344]==1) 
	 		intermediate[4095+2344:0+2344] <= intermediate[4095+2344:0+2344] + a; end
12'd2345: begin if(a[2345]==1) 
	 		intermediate[4095+2345:0+2345] <= intermediate[4095+2345:0+2345] + a; end
12'd2346: begin if(a[2346]==1) 
	 		intermediate[4095+2346:0+2346] <= intermediate[4095+2346:0+2346] + a; end
12'd2347: begin if(a[2347]==1) 
	 		intermediate[4095+2347:0+2347] <= intermediate[4095+2347:0+2347] + a; end
12'd2348: begin if(a[2348]==1) 
	 		intermediate[4095+2348:0+2348] <= intermediate[4095+2348:0+2348] + a; end
12'd2349: begin if(a[2349]==1) 
	 		intermediate[4095+2349:0+2349] <= intermediate[4095+2349:0+2349] + a; end
12'd2350: begin if(a[2350]==1) 
	 		intermediate[4095+2350:0+2350] <= intermediate[4095+2350:0+2350] + a; end
12'd2351: begin if(a[2351]==1) 
	 		intermediate[4095+2351:0+2351] <= intermediate[4095+2351:0+2351] + a; end
12'd2352: begin if(a[2352]==1) 
	 		intermediate[4095+2352:0+2352] <= intermediate[4095+2352:0+2352] + a; end
12'd2353: begin if(a[2353]==1) 
	 		intermediate[4095+2353:0+2353] <= intermediate[4095+2353:0+2353] + a; end
12'd2354: begin if(a[2354]==1) 
	 		intermediate[4095+2354:0+2354] <= intermediate[4095+2354:0+2354] + a; end
12'd2355: begin if(a[2355]==1) 
	 		intermediate[4095+2355:0+2355] <= intermediate[4095+2355:0+2355] + a; end
12'd2356: begin if(a[2356]==1) 
	 		intermediate[4095+2356:0+2356] <= intermediate[4095+2356:0+2356] + a; end
12'd2357: begin if(a[2357]==1) 
	 		intermediate[4095+2357:0+2357] <= intermediate[4095+2357:0+2357] + a; end
12'd2358: begin if(a[2358]==1) 
	 		intermediate[4095+2358:0+2358] <= intermediate[4095+2358:0+2358] + a; end
12'd2359: begin if(a[2359]==1) 
	 		intermediate[4095+2359:0+2359] <= intermediate[4095+2359:0+2359] + a; end
12'd2360: begin if(a[2360]==1) 
	 		intermediate[4095+2360:0+2360] <= intermediate[4095+2360:0+2360] + a; end
12'd2361: begin if(a[2361]==1) 
	 		intermediate[4095+2361:0+2361] <= intermediate[4095+2361:0+2361] + a; end
12'd2362: begin if(a[2362]==1) 
	 		intermediate[4095+2362:0+2362] <= intermediate[4095+2362:0+2362] + a; end
12'd2363: begin if(a[2363]==1) 
	 		intermediate[4095+2363:0+2363] <= intermediate[4095+2363:0+2363] + a; end
12'd2364: begin if(a[2364]==1) 
	 		intermediate[4095+2364:0+2364] <= intermediate[4095+2364:0+2364] + a; end
12'd2365: begin if(a[2365]==1) 
	 		intermediate[4095+2365:0+2365] <= intermediate[4095+2365:0+2365] + a; end
12'd2366: begin if(a[2366]==1) 
	 		intermediate[4095+2366:0+2366] <= intermediate[4095+2366:0+2366] + a; end
12'd2367: begin if(a[2367]==1) 
	 		intermediate[4095+2367:0+2367] <= intermediate[4095+2367:0+2367] + a; end
12'd2368: begin if(a[2368]==1) 
	 		intermediate[4095+2368:0+2368] <= intermediate[4095+2368:0+2368] + a; end
12'd2369: begin if(a[2369]==1) 
	 		intermediate[4095+2369:0+2369] <= intermediate[4095+2369:0+2369] + a; end
12'd2370: begin if(a[2370]==1) 
	 		intermediate[4095+2370:0+2370] <= intermediate[4095+2370:0+2370] + a; end
12'd2371: begin if(a[2371]==1) 
	 		intermediate[4095+2371:0+2371] <= intermediate[4095+2371:0+2371] + a; end
12'd2372: begin if(a[2372]==1) 
	 		intermediate[4095+2372:0+2372] <= intermediate[4095+2372:0+2372] + a; end
12'd2373: begin if(a[2373]==1) 
	 		intermediate[4095+2373:0+2373] <= intermediate[4095+2373:0+2373] + a; end
12'd2374: begin if(a[2374]==1) 
	 		intermediate[4095+2374:0+2374] <= intermediate[4095+2374:0+2374] + a; end
12'd2375: begin if(a[2375]==1) 
	 		intermediate[4095+2375:0+2375] <= intermediate[4095+2375:0+2375] + a; end
12'd2376: begin if(a[2376]==1) 
	 		intermediate[4095+2376:0+2376] <= intermediate[4095+2376:0+2376] + a; end
12'd2377: begin if(a[2377]==1) 
	 		intermediate[4095+2377:0+2377] <= intermediate[4095+2377:0+2377] + a; end
12'd2378: begin if(a[2378]==1) 
	 		intermediate[4095+2378:0+2378] <= intermediate[4095+2378:0+2378] + a; end
12'd2379: begin if(a[2379]==1) 
	 		intermediate[4095+2379:0+2379] <= intermediate[4095+2379:0+2379] + a; end
12'd2380: begin if(a[2380]==1) 
	 		intermediate[4095+2380:0+2380] <= intermediate[4095+2380:0+2380] + a; end
12'd2381: begin if(a[2381]==1) 
	 		intermediate[4095+2381:0+2381] <= intermediate[4095+2381:0+2381] + a; end
12'd2382: begin if(a[2382]==1) 
	 		intermediate[4095+2382:0+2382] <= intermediate[4095+2382:0+2382] + a; end
12'd2383: begin if(a[2383]==1) 
	 		intermediate[4095+2383:0+2383] <= intermediate[4095+2383:0+2383] + a; end
12'd2384: begin if(a[2384]==1) 
	 		intermediate[4095+2384:0+2384] <= intermediate[4095+2384:0+2384] + a; end
12'd2385: begin if(a[2385]==1) 
	 		intermediate[4095+2385:0+2385] <= intermediate[4095+2385:0+2385] + a; end
12'd2386: begin if(a[2386]==1) 
	 		intermediate[4095+2386:0+2386] <= intermediate[4095+2386:0+2386] + a; end
12'd2387: begin if(a[2387]==1) 
	 		intermediate[4095+2387:0+2387] <= intermediate[4095+2387:0+2387] + a; end
12'd2388: begin if(a[2388]==1) 
	 		intermediate[4095+2388:0+2388] <= intermediate[4095+2388:0+2388] + a; end
12'd2389: begin if(a[2389]==1) 
	 		intermediate[4095+2389:0+2389] <= intermediate[4095+2389:0+2389] + a; end
12'd2390: begin if(a[2390]==1) 
	 		intermediate[4095+2390:0+2390] <= intermediate[4095+2390:0+2390] + a; end
12'd2391: begin if(a[2391]==1) 
	 		intermediate[4095+2391:0+2391] <= intermediate[4095+2391:0+2391] + a; end
12'd2392: begin if(a[2392]==1) 
	 		intermediate[4095+2392:0+2392] <= intermediate[4095+2392:0+2392] + a; end
12'd2393: begin if(a[2393]==1) 
	 		intermediate[4095+2393:0+2393] <= intermediate[4095+2393:0+2393] + a; end
12'd2394: begin if(a[2394]==1) 
	 		intermediate[4095+2394:0+2394] <= intermediate[4095+2394:0+2394] + a; end
12'd2395: begin if(a[2395]==1) 
	 		intermediate[4095+2395:0+2395] <= intermediate[4095+2395:0+2395] + a; end
12'd2396: begin if(a[2396]==1) 
	 		intermediate[4095+2396:0+2396] <= intermediate[4095+2396:0+2396] + a; end
12'd2397: begin if(a[2397]==1) 
	 		intermediate[4095+2397:0+2397] <= intermediate[4095+2397:0+2397] + a; end
12'd2398: begin if(a[2398]==1) 
	 		intermediate[4095+2398:0+2398] <= intermediate[4095+2398:0+2398] + a; end
12'd2399: begin if(a[2399]==1) 
	 		intermediate[4095+2399:0+2399] <= intermediate[4095+2399:0+2399] + a; end
12'd2400: begin if(a[2400]==1) 
	 		intermediate[4095+2400:0+2400] <= intermediate[4095+2400:0+2400] + a; end
12'd2401: begin if(a[2401]==1) 
	 		intermediate[4095+2401:0+2401] <= intermediate[4095+2401:0+2401] + a; end
12'd2402: begin if(a[2402]==1) 
	 		intermediate[4095+2402:0+2402] <= intermediate[4095+2402:0+2402] + a; end
12'd2403: begin if(a[2403]==1) 
	 		intermediate[4095+2403:0+2403] <= intermediate[4095+2403:0+2403] + a; end
12'd2404: begin if(a[2404]==1) 
	 		intermediate[4095+2404:0+2404] <= intermediate[4095+2404:0+2404] + a; end
12'd2405: begin if(a[2405]==1) 
	 		intermediate[4095+2405:0+2405] <= intermediate[4095+2405:0+2405] + a; end
12'd2406: begin if(a[2406]==1) 
	 		intermediate[4095+2406:0+2406] <= intermediate[4095+2406:0+2406] + a; end
12'd2407: begin if(a[2407]==1) 
	 		intermediate[4095+2407:0+2407] <= intermediate[4095+2407:0+2407] + a; end
12'd2408: begin if(a[2408]==1) 
	 		intermediate[4095+2408:0+2408] <= intermediate[4095+2408:0+2408] + a; end
12'd2409: begin if(a[2409]==1) 
	 		intermediate[4095+2409:0+2409] <= intermediate[4095+2409:0+2409] + a; end
12'd2410: begin if(a[2410]==1) 
	 		intermediate[4095+2410:0+2410] <= intermediate[4095+2410:0+2410] + a; end
12'd2411: begin if(a[2411]==1) 
	 		intermediate[4095+2411:0+2411] <= intermediate[4095+2411:0+2411] + a; end
12'd2412: begin if(a[2412]==1) 
	 		intermediate[4095+2412:0+2412] <= intermediate[4095+2412:0+2412] + a; end
12'd2413: begin if(a[2413]==1) 
	 		intermediate[4095+2413:0+2413] <= intermediate[4095+2413:0+2413] + a; end
12'd2414: begin if(a[2414]==1) 
	 		intermediate[4095+2414:0+2414] <= intermediate[4095+2414:0+2414] + a; end
12'd2415: begin if(a[2415]==1) 
	 		intermediate[4095+2415:0+2415] <= intermediate[4095+2415:0+2415] + a; end
12'd2416: begin if(a[2416]==1) 
	 		intermediate[4095+2416:0+2416] <= intermediate[4095+2416:0+2416] + a; end
12'd2417: begin if(a[2417]==1) 
	 		intermediate[4095+2417:0+2417] <= intermediate[4095+2417:0+2417] + a; end
12'd2418: begin if(a[2418]==1) 
	 		intermediate[4095+2418:0+2418] <= intermediate[4095+2418:0+2418] + a; end
12'd2419: begin if(a[2419]==1) 
	 		intermediate[4095+2419:0+2419] <= intermediate[4095+2419:0+2419] + a; end
12'd2420: begin if(a[2420]==1) 
	 		intermediate[4095+2420:0+2420] <= intermediate[4095+2420:0+2420] + a; end
12'd2421: begin if(a[2421]==1) 
	 		intermediate[4095+2421:0+2421] <= intermediate[4095+2421:0+2421] + a; end
12'd2422: begin if(a[2422]==1) 
	 		intermediate[4095+2422:0+2422] <= intermediate[4095+2422:0+2422] + a; end
12'd2423: begin if(a[2423]==1) 
	 		intermediate[4095+2423:0+2423] <= intermediate[4095+2423:0+2423] + a; end
12'd2424: begin if(a[2424]==1) 
	 		intermediate[4095+2424:0+2424] <= intermediate[4095+2424:0+2424] + a; end
12'd2425: begin if(a[2425]==1) 
	 		intermediate[4095+2425:0+2425] <= intermediate[4095+2425:0+2425] + a; end
12'd2426: begin if(a[2426]==1) 
	 		intermediate[4095+2426:0+2426] <= intermediate[4095+2426:0+2426] + a; end
12'd2427: begin if(a[2427]==1) 
	 		intermediate[4095+2427:0+2427] <= intermediate[4095+2427:0+2427] + a; end
12'd2428: begin if(a[2428]==1) 
	 		intermediate[4095+2428:0+2428] <= intermediate[4095+2428:0+2428] + a; end
12'd2429: begin if(a[2429]==1) 
	 		intermediate[4095+2429:0+2429] <= intermediate[4095+2429:0+2429] + a; end
12'd2430: begin if(a[2430]==1) 
	 		intermediate[4095+2430:0+2430] <= intermediate[4095+2430:0+2430] + a; end
12'd2431: begin if(a[2431]==1) 
	 		intermediate[4095+2431:0+2431] <= intermediate[4095+2431:0+2431] + a; end
12'd2432: begin if(a[2432]==1) 
	 		intermediate[4095+2432:0+2432] <= intermediate[4095+2432:0+2432] + a; end
12'd2433: begin if(a[2433]==1) 
	 		intermediate[4095+2433:0+2433] <= intermediate[4095+2433:0+2433] + a; end
12'd2434: begin if(a[2434]==1) 
	 		intermediate[4095+2434:0+2434] <= intermediate[4095+2434:0+2434] + a; end
12'd2435: begin if(a[2435]==1) 
	 		intermediate[4095+2435:0+2435] <= intermediate[4095+2435:0+2435] + a; end
12'd2436: begin if(a[2436]==1) 
	 		intermediate[4095+2436:0+2436] <= intermediate[4095+2436:0+2436] + a; end
12'd2437: begin if(a[2437]==1) 
	 		intermediate[4095+2437:0+2437] <= intermediate[4095+2437:0+2437] + a; end
12'd2438: begin if(a[2438]==1) 
	 		intermediate[4095+2438:0+2438] <= intermediate[4095+2438:0+2438] + a; end
12'd2439: begin if(a[2439]==1) 
	 		intermediate[4095+2439:0+2439] <= intermediate[4095+2439:0+2439] + a; end
12'd2440: begin if(a[2440]==1) 
	 		intermediate[4095+2440:0+2440] <= intermediate[4095+2440:0+2440] + a; end
12'd2441: begin if(a[2441]==1) 
	 		intermediate[4095+2441:0+2441] <= intermediate[4095+2441:0+2441] + a; end
12'd2442: begin if(a[2442]==1) 
	 		intermediate[4095+2442:0+2442] <= intermediate[4095+2442:0+2442] + a; end
12'd2443: begin if(a[2443]==1) 
	 		intermediate[4095+2443:0+2443] <= intermediate[4095+2443:0+2443] + a; end
12'd2444: begin if(a[2444]==1) 
	 		intermediate[4095+2444:0+2444] <= intermediate[4095+2444:0+2444] + a; end
12'd2445: begin if(a[2445]==1) 
	 		intermediate[4095+2445:0+2445] <= intermediate[4095+2445:0+2445] + a; end
12'd2446: begin if(a[2446]==1) 
	 		intermediate[4095+2446:0+2446] <= intermediate[4095+2446:0+2446] + a; end
12'd2447: begin if(a[2447]==1) 
	 		intermediate[4095+2447:0+2447] <= intermediate[4095+2447:0+2447] + a; end
12'd2448: begin if(a[2448]==1) 
	 		intermediate[4095+2448:0+2448] <= intermediate[4095+2448:0+2448] + a; end
12'd2449: begin if(a[2449]==1) 
	 		intermediate[4095+2449:0+2449] <= intermediate[4095+2449:0+2449] + a; end
12'd2450: begin if(a[2450]==1) 
	 		intermediate[4095+2450:0+2450] <= intermediate[4095+2450:0+2450] + a; end
12'd2451: begin if(a[2451]==1) 
	 		intermediate[4095+2451:0+2451] <= intermediate[4095+2451:0+2451] + a; end
12'd2452: begin if(a[2452]==1) 
	 		intermediate[4095+2452:0+2452] <= intermediate[4095+2452:0+2452] + a; end
12'd2453: begin if(a[2453]==1) 
	 		intermediate[4095+2453:0+2453] <= intermediate[4095+2453:0+2453] + a; end
12'd2454: begin if(a[2454]==1) 
	 		intermediate[4095+2454:0+2454] <= intermediate[4095+2454:0+2454] + a; end
12'd2455: begin if(a[2455]==1) 
	 		intermediate[4095+2455:0+2455] <= intermediate[4095+2455:0+2455] + a; end
12'd2456: begin if(a[2456]==1) 
	 		intermediate[4095+2456:0+2456] <= intermediate[4095+2456:0+2456] + a; end
12'd2457: begin if(a[2457]==1) 
	 		intermediate[4095+2457:0+2457] <= intermediate[4095+2457:0+2457] + a; end
12'd2458: begin if(a[2458]==1) 
	 		intermediate[4095+2458:0+2458] <= intermediate[4095+2458:0+2458] + a; end
12'd2459: begin if(a[2459]==1) 
	 		intermediate[4095+2459:0+2459] <= intermediate[4095+2459:0+2459] + a; end
12'd2460: begin if(a[2460]==1) 
	 		intermediate[4095+2460:0+2460] <= intermediate[4095+2460:0+2460] + a; end
12'd2461: begin if(a[2461]==1) 
	 		intermediate[4095+2461:0+2461] <= intermediate[4095+2461:0+2461] + a; end
12'd2462: begin if(a[2462]==1) 
	 		intermediate[4095+2462:0+2462] <= intermediate[4095+2462:0+2462] + a; end
12'd2463: begin if(a[2463]==1) 
	 		intermediate[4095+2463:0+2463] <= intermediate[4095+2463:0+2463] + a; end
12'd2464: begin if(a[2464]==1) 
	 		intermediate[4095+2464:0+2464] <= intermediate[4095+2464:0+2464] + a; end
12'd2465: begin if(a[2465]==1) 
	 		intermediate[4095+2465:0+2465] <= intermediate[4095+2465:0+2465] + a; end
12'd2466: begin if(a[2466]==1) 
	 		intermediate[4095+2466:0+2466] <= intermediate[4095+2466:0+2466] + a; end
12'd2467: begin if(a[2467]==1) 
	 		intermediate[4095+2467:0+2467] <= intermediate[4095+2467:0+2467] + a; end
12'd2468: begin if(a[2468]==1) 
	 		intermediate[4095+2468:0+2468] <= intermediate[4095+2468:0+2468] + a; end
12'd2469: begin if(a[2469]==1) 
	 		intermediate[4095+2469:0+2469] <= intermediate[4095+2469:0+2469] + a; end
12'd2470: begin if(a[2470]==1) 
	 		intermediate[4095+2470:0+2470] <= intermediate[4095+2470:0+2470] + a; end
12'd2471: begin if(a[2471]==1) 
	 		intermediate[4095+2471:0+2471] <= intermediate[4095+2471:0+2471] + a; end
12'd2472: begin if(a[2472]==1) 
	 		intermediate[4095+2472:0+2472] <= intermediate[4095+2472:0+2472] + a; end
12'd2473: begin if(a[2473]==1) 
	 		intermediate[4095+2473:0+2473] <= intermediate[4095+2473:0+2473] + a; end
12'd2474: begin if(a[2474]==1) 
	 		intermediate[4095+2474:0+2474] <= intermediate[4095+2474:0+2474] + a; end
12'd2475: begin if(a[2475]==1) 
	 		intermediate[4095+2475:0+2475] <= intermediate[4095+2475:0+2475] + a; end
12'd2476: begin if(a[2476]==1) 
	 		intermediate[4095+2476:0+2476] <= intermediate[4095+2476:0+2476] + a; end
12'd2477: begin if(a[2477]==1) 
	 		intermediate[4095+2477:0+2477] <= intermediate[4095+2477:0+2477] + a; end
12'd2478: begin if(a[2478]==1) 
	 		intermediate[4095+2478:0+2478] <= intermediate[4095+2478:0+2478] + a; end
12'd2479: begin if(a[2479]==1) 
	 		intermediate[4095+2479:0+2479] <= intermediate[4095+2479:0+2479] + a; end
12'd2480: begin if(a[2480]==1) 
	 		intermediate[4095+2480:0+2480] <= intermediate[4095+2480:0+2480] + a; end
12'd2481: begin if(a[2481]==1) 
	 		intermediate[4095+2481:0+2481] <= intermediate[4095+2481:0+2481] + a; end
12'd2482: begin if(a[2482]==1) 
	 		intermediate[4095+2482:0+2482] <= intermediate[4095+2482:0+2482] + a; end
12'd2483: begin if(a[2483]==1) 
	 		intermediate[4095+2483:0+2483] <= intermediate[4095+2483:0+2483] + a; end
12'd2484: begin if(a[2484]==1) 
	 		intermediate[4095+2484:0+2484] <= intermediate[4095+2484:0+2484] + a; end
12'd2485: begin if(a[2485]==1) 
	 		intermediate[4095+2485:0+2485] <= intermediate[4095+2485:0+2485] + a; end
12'd2486: begin if(a[2486]==1) 
	 		intermediate[4095+2486:0+2486] <= intermediate[4095+2486:0+2486] + a; end
12'd2487: begin if(a[2487]==1) 
	 		intermediate[4095+2487:0+2487] <= intermediate[4095+2487:0+2487] + a; end
12'd2488: begin if(a[2488]==1) 
	 		intermediate[4095+2488:0+2488] <= intermediate[4095+2488:0+2488] + a; end
12'd2489: begin if(a[2489]==1) 
	 		intermediate[4095+2489:0+2489] <= intermediate[4095+2489:0+2489] + a; end
12'd2490: begin if(a[2490]==1) 
	 		intermediate[4095+2490:0+2490] <= intermediate[4095+2490:0+2490] + a; end
12'd2491: begin if(a[2491]==1) 
	 		intermediate[4095+2491:0+2491] <= intermediate[4095+2491:0+2491] + a; end
12'd2492: begin if(a[2492]==1) 
	 		intermediate[4095+2492:0+2492] <= intermediate[4095+2492:0+2492] + a; end
12'd2493: begin if(a[2493]==1) 
	 		intermediate[4095+2493:0+2493] <= intermediate[4095+2493:0+2493] + a; end
12'd2494: begin if(a[2494]==1) 
	 		intermediate[4095+2494:0+2494] <= intermediate[4095+2494:0+2494] + a; end
12'd2495: begin if(a[2495]==1) 
	 		intermediate[4095+2495:0+2495] <= intermediate[4095+2495:0+2495] + a; end
12'd2496: begin if(a[2496]==1) 
	 		intermediate[4095+2496:0+2496] <= intermediate[4095+2496:0+2496] + a; end
12'd2497: begin if(a[2497]==1) 
	 		intermediate[4095+2497:0+2497] <= intermediate[4095+2497:0+2497] + a; end
12'd2498: begin if(a[2498]==1) 
	 		intermediate[4095+2498:0+2498] <= intermediate[4095+2498:0+2498] + a; end
12'd2499: begin if(a[2499]==1) 
	 		intermediate[4095+2499:0+2499] <= intermediate[4095+2499:0+2499] + a; end
12'd2500: begin if(a[2500]==1) 
	 		intermediate[4095+2500:0+2500] <= intermediate[4095+2500:0+2500] + a; end
12'd2501: begin if(a[2501]==1) 
	 		intermediate[4095+2501:0+2501] <= intermediate[4095+2501:0+2501] + a; end
12'd2502: begin if(a[2502]==1) 
	 		intermediate[4095+2502:0+2502] <= intermediate[4095+2502:0+2502] + a; end
12'd2503: begin if(a[2503]==1) 
	 		intermediate[4095+2503:0+2503] <= intermediate[4095+2503:0+2503] + a; end
12'd2504: begin if(a[2504]==1) 
	 		intermediate[4095+2504:0+2504] <= intermediate[4095+2504:0+2504] + a; end
12'd2505: begin if(a[2505]==1) 
	 		intermediate[4095+2505:0+2505] <= intermediate[4095+2505:0+2505] + a; end
12'd2506: begin if(a[2506]==1) 
	 		intermediate[4095+2506:0+2506] <= intermediate[4095+2506:0+2506] + a; end
12'd2507: begin if(a[2507]==1) 
	 		intermediate[4095+2507:0+2507] <= intermediate[4095+2507:0+2507] + a; end
12'd2508: begin if(a[2508]==1) 
	 		intermediate[4095+2508:0+2508] <= intermediate[4095+2508:0+2508] + a; end
12'd2509: begin if(a[2509]==1) 
	 		intermediate[4095+2509:0+2509] <= intermediate[4095+2509:0+2509] + a; end
12'd2510: begin if(a[2510]==1) 
	 		intermediate[4095+2510:0+2510] <= intermediate[4095+2510:0+2510] + a; end
12'd2511: begin if(a[2511]==1) 
	 		intermediate[4095+2511:0+2511] <= intermediate[4095+2511:0+2511] + a; end
12'd2512: begin if(a[2512]==1) 
	 		intermediate[4095+2512:0+2512] <= intermediate[4095+2512:0+2512] + a; end
12'd2513: begin if(a[2513]==1) 
	 		intermediate[4095+2513:0+2513] <= intermediate[4095+2513:0+2513] + a; end
12'd2514: begin if(a[2514]==1) 
	 		intermediate[4095+2514:0+2514] <= intermediate[4095+2514:0+2514] + a; end
12'd2515: begin if(a[2515]==1) 
	 		intermediate[4095+2515:0+2515] <= intermediate[4095+2515:0+2515] + a; end
12'd2516: begin if(a[2516]==1) 
	 		intermediate[4095+2516:0+2516] <= intermediate[4095+2516:0+2516] + a; end
12'd2517: begin if(a[2517]==1) 
	 		intermediate[4095+2517:0+2517] <= intermediate[4095+2517:0+2517] + a; end
12'd2518: begin if(a[2518]==1) 
	 		intermediate[4095+2518:0+2518] <= intermediate[4095+2518:0+2518] + a; end
12'd2519: begin if(a[2519]==1) 
	 		intermediate[4095+2519:0+2519] <= intermediate[4095+2519:0+2519] + a; end
12'd2520: begin if(a[2520]==1) 
	 		intermediate[4095+2520:0+2520] <= intermediate[4095+2520:0+2520] + a; end
12'd2521: begin if(a[2521]==1) 
	 		intermediate[4095+2521:0+2521] <= intermediate[4095+2521:0+2521] + a; end
12'd2522: begin if(a[2522]==1) 
	 		intermediate[4095+2522:0+2522] <= intermediate[4095+2522:0+2522] + a; end
12'd2523: begin if(a[2523]==1) 
	 		intermediate[4095+2523:0+2523] <= intermediate[4095+2523:0+2523] + a; end
12'd2524: begin if(a[2524]==1) 
	 		intermediate[4095+2524:0+2524] <= intermediate[4095+2524:0+2524] + a; end
12'd2525: begin if(a[2525]==1) 
	 		intermediate[4095+2525:0+2525] <= intermediate[4095+2525:0+2525] + a; end
12'd2526: begin if(a[2526]==1) 
	 		intermediate[4095+2526:0+2526] <= intermediate[4095+2526:0+2526] + a; end
12'd2527: begin if(a[2527]==1) 
	 		intermediate[4095+2527:0+2527] <= intermediate[4095+2527:0+2527] + a; end
12'd2528: begin if(a[2528]==1) 
	 		intermediate[4095+2528:0+2528] <= intermediate[4095+2528:0+2528] + a; end
12'd2529: begin if(a[2529]==1) 
	 		intermediate[4095+2529:0+2529] <= intermediate[4095+2529:0+2529] + a; end
12'd2530: begin if(a[2530]==1) 
	 		intermediate[4095+2530:0+2530] <= intermediate[4095+2530:0+2530] + a; end
12'd2531: begin if(a[2531]==1) 
	 		intermediate[4095+2531:0+2531] <= intermediate[4095+2531:0+2531] + a; end
12'd2532: begin if(a[2532]==1) 
	 		intermediate[4095+2532:0+2532] <= intermediate[4095+2532:0+2532] + a; end
12'd2533: begin if(a[2533]==1) 
	 		intermediate[4095+2533:0+2533] <= intermediate[4095+2533:0+2533] + a; end
12'd2534: begin if(a[2534]==1) 
	 		intermediate[4095+2534:0+2534] <= intermediate[4095+2534:0+2534] + a; end
12'd2535: begin if(a[2535]==1) 
	 		intermediate[4095+2535:0+2535] <= intermediate[4095+2535:0+2535] + a; end
12'd2536: begin if(a[2536]==1) 
	 		intermediate[4095+2536:0+2536] <= intermediate[4095+2536:0+2536] + a; end
12'd2537: begin if(a[2537]==1) 
	 		intermediate[4095+2537:0+2537] <= intermediate[4095+2537:0+2537] + a; end
12'd2538: begin if(a[2538]==1) 
	 		intermediate[4095+2538:0+2538] <= intermediate[4095+2538:0+2538] + a; end
12'd2539: begin if(a[2539]==1) 
	 		intermediate[4095+2539:0+2539] <= intermediate[4095+2539:0+2539] + a; end
12'd2540: begin if(a[2540]==1) 
	 		intermediate[4095+2540:0+2540] <= intermediate[4095+2540:0+2540] + a; end
12'd2541: begin if(a[2541]==1) 
	 		intermediate[4095+2541:0+2541] <= intermediate[4095+2541:0+2541] + a; end
12'd2542: begin if(a[2542]==1) 
	 		intermediate[4095+2542:0+2542] <= intermediate[4095+2542:0+2542] + a; end
12'd2543: begin if(a[2543]==1) 
	 		intermediate[4095+2543:0+2543] <= intermediate[4095+2543:0+2543] + a; end
12'd2544: begin if(a[2544]==1) 
	 		intermediate[4095+2544:0+2544] <= intermediate[4095+2544:0+2544] + a; end
12'd2545: begin if(a[2545]==1) 
	 		intermediate[4095+2545:0+2545] <= intermediate[4095+2545:0+2545] + a; end
12'd2546: begin if(a[2546]==1) 
	 		intermediate[4095+2546:0+2546] <= intermediate[4095+2546:0+2546] + a; end
12'd2547: begin if(a[2547]==1) 
	 		intermediate[4095+2547:0+2547] <= intermediate[4095+2547:0+2547] + a; end
12'd2548: begin if(a[2548]==1) 
	 		intermediate[4095+2548:0+2548] <= intermediate[4095+2548:0+2548] + a; end
12'd2549: begin if(a[2549]==1) 
	 		intermediate[4095+2549:0+2549] <= intermediate[4095+2549:0+2549] + a; end
12'd2550: begin if(a[2550]==1) 
	 		intermediate[4095+2550:0+2550] <= intermediate[4095+2550:0+2550] + a; end
12'd2551: begin if(a[2551]==1) 
	 		intermediate[4095+2551:0+2551] <= intermediate[4095+2551:0+2551] + a; end
12'd2552: begin if(a[2552]==1) 
	 		intermediate[4095+2552:0+2552] <= intermediate[4095+2552:0+2552] + a; end
12'd2553: begin if(a[2553]==1) 
	 		intermediate[4095+2553:0+2553] <= intermediate[4095+2553:0+2553] + a; end
12'd2554: begin if(a[2554]==1) 
	 		intermediate[4095+2554:0+2554] <= intermediate[4095+2554:0+2554] + a; end
12'd2555: begin if(a[2555]==1) 
	 		intermediate[4095+2555:0+2555] <= intermediate[4095+2555:0+2555] + a; end
12'd2556: begin if(a[2556]==1) 
	 		intermediate[4095+2556:0+2556] <= intermediate[4095+2556:0+2556] + a; end
12'd2557: begin if(a[2557]==1) 
	 		intermediate[4095+2557:0+2557] <= intermediate[4095+2557:0+2557] + a; end
12'd2558: begin if(a[2558]==1) 
	 		intermediate[4095+2558:0+2558] <= intermediate[4095+2558:0+2558] + a; end
12'd2559: begin if(a[2559]==1) 
	 		intermediate[4095+2559:0+2559] <= intermediate[4095+2559:0+2559] + a; end
12'd2560: begin if(a[2560]==1) 
	 		intermediate[4095+2560:0+2560] <= intermediate[4095+2560:0+2560] + a; end
12'd2561: begin if(a[2561]==1) 
	 		intermediate[4095+2561:0+2561] <= intermediate[4095+2561:0+2561] + a; end
12'd2562: begin if(a[2562]==1) 
	 		intermediate[4095+2562:0+2562] <= intermediate[4095+2562:0+2562] + a; end
12'd2563: begin if(a[2563]==1) 
	 		intermediate[4095+2563:0+2563] <= intermediate[4095+2563:0+2563] + a; end
12'd2564: begin if(a[2564]==1) 
	 		intermediate[4095+2564:0+2564] <= intermediate[4095+2564:0+2564] + a; end
12'd2565: begin if(a[2565]==1) 
	 		intermediate[4095+2565:0+2565] <= intermediate[4095+2565:0+2565] + a; end
12'd2566: begin if(a[2566]==1) 
	 		intermediate[4095+2566:0+2566] <= intermediate[4095+2566:0+2566] + a; end
12'd2567: begin if(a[2567]==1) 
	 		intermediate[4095+2567:0+2567] <= intermediate[4095+2567:0+2567] + a; end
12'd2568: begin if(a[2568]==1) 
	 		intermediate[4095+2568:0+2568] <= intermediate[4095+2568:0+2568] + a; end
12'd2569: begin if(a[2569]==1) 
	 		intermediate[4095+2569:0+2569] <= intermediate[4095+2569:0+2569] + a; end
12'd2570: begin if(a[2570]==1) 
	 		intermediate[4095+2570:0+2570] <= intermediate[4095+2570:0+2570] + a; end
12'd2571: begin if(a[2571]==1) 
	 		intermediate[4095+2571:0+2571] <= intermediate[4095+2571:0+2571] + a; end
12'd2572: begin if(a[2572]==1) 
	 		intermediate[4095+2572:0+2572] <= intermediate[4095+2572:0+2572] + a; end
12'd2573: begin if(a[2573]==1) 
	 		intermediate[4095+2573:0+2573] <= intermediate[4095+2573:0+2573] + a; end
12'd2574: begin if(a[2574]==1) 
	 		intermediate[4095+2574:0+2574] <= intermediate[4095+2574:0+2574] + a; end
12'd2575: begin if(a[2575]==1) 
	 		intermediate[4095+2575:0+2575] <= intermediate[4095+2575:0+2575] + a; end
12'd2576: begin if(a[2576]==1) 
	 		intermediate[4095+2576:0+2576] <= intermediate[4095+2576:0+2576] + a; end
12'd2577: begin if(a[2577]==1) 
	 		intermediate[4095+2577:0+2577] <= intermediate[4095+2577:0+2577] + a; end
12'd2578: begin if(a[2578]==1) 
	 		intermediate[4095+2578:0+2578] <= intermediate[4095+2578:0+2578] + a; end
12'd2579: begin if(a[2579]==1) 
	 		intermediate[4095+2579:0+2579] <= intermediate[4095+2579:0+2579] + a; end
12'd2580: begin if(a[2580]==1) 
	 		intermediate[4095+2580:0+2580] <= intermediate[4095+2580:0+2580] + a; end
12'd2581: begin if(a[2581]==1) 
	 		intermediate[4095+2581:0+2581] <= intermediate[4095+2581:0+2581] + a; end
12'd2582: begin if(a[2582]==1) 
	 		intermediate[4095+2582:0+2582] <= intermediate[4095+2582:0+2582] + a; end
12'd2583: begin if(a[2583]==1) 
	 		intermediate[4095+2583:0+2583] <= intermediate[4095+2583:0+2583] + a; end
12'd2584: begin if(a[2584]==1) 
	 		intermediate[4095+2584:0+2584] <= intermediate[4095+2584:0+2584] + a; end
12'd2585: begin if(a[2585]==1) 
	 		intermediate[4095+2585:0+2585] <= intermediate[4095+2585:0+2585] + a; end
12'd2586: begin if(a[2586]==1) 
	 		intermediate[4095+2586:0+2586] <= intermediate[4095+2586:0+2586] + a; end
12'd2587: begin if(a[2587]==1) 
	 		intermediate[4095+2587:0+2587] <= intermediate[4095+2587:0+2587] + a; end
12'd2588: begin if(a[2588]==1) 
	 		intermediate[4095+2588:0+2588] <= intermediate[4095+2588:0+2588] + a; end
12'd2589: begin if(a[2589]==1) 
	 		intermediate[4095+2589:0+2589] <= intermediate[4095+2589:0+2589] + a; end
12'd2590: begin if(a[2590]==1) 
	 		intermediate[4095+2590:0+2590] <= intermediate[4095+2590:0+2590] + a; end
12'd2591: begin if(a[2591]==1) 
	 		intermediate[4095+2591:0+2591] <= intermediate[4095+2591:0+2591] + a; end
12'd2592: begin if(a[2592]==1) 
	 		intermediate[4095+2592:0+2592] <= intermediate[4095+2592:0+2592] + a; end
12'd2593: begin if(a[2593]==1) 
	 		intermediate[4095+2593:0+2593] <= intermediate[4095+2593:0+2593] + a; end
12'd2594: begin if(a[2594]==1) 
	 		intermediate[4095+2594:0+2594] <= intermediate[4095+2594:0+2594] + a; end
12'd2595: begin if(a[2595]==1) 
	 		intermediate[4095+2595:0+2595] <= intermediate[4095+2595:0+2595] + a; end
12'd2596: begin if(a[2596]==1) 
	 		intermediate[4095+2596:0+2596] <= intermediate[4095+2596:0+2596] + a; end
12'd2597: begin if(a[2597]==1) 
	 		intermediate[4095+2597:0+2597] <= intermediate[4095+2597:0+2597] + a; end
12'd2598: begin if(a[2598]==1) 
	 		intermediate[4095+2598:0+2598] <= intermediate[4095+2598:0+2598] + a; end
12'd2599: begin if(a[2599]==1) 
	 		intermediate[4095+2599:0+2599] <= intermediate[4095+2599:0+2599] + a; end
12'd2600: begin if(a[2600]==1) 
	 		intermediate[4095+2600:0+2600] <= intermediate[4095+2600:0+2600] + a; end
12'd2601: begin if(a[2601]==1) 
	 		intermediate[4095+2601:0+2601] <= intermediate[4095+2601:0+2601] + a; end
12'd2602: begin if(a[2602]==1) 
	 		intermediate[4095+2602:0+2602] <= intermediate[4095+2602:0+2602] + a; end
12'd2603: begin if(a[2603]==1) 
	 		intermediate[4095+2603:0+2603] <= intermediate[4095+2603:0+2603] + a; end
12'd2604: begin if(a[2604]==1) 
	 		intermediate[4095+2604:0+2604] <= intermediate[4095+2604:0+2604] + a; end
12'd2605: begin if(a[2605]==1) 
	 		intermediate[4095+2605:0+2605] <= intermediate[4095+2605:0+2605] + a; end
12'd2606: begin if(a[2606]==1) 
	 		intermediate[4095+2606:0+2606] <= intermediate[4095+2606:0+2606] + a; end
12'd2607: begin if(a[2607]==1) 
	 		intermediate[4095+2607:0+2607] <= intermediate[4095+2607:0+2607] + a; end
12'd2608: begin if(a[2608]==1) 
	 		intermediate[4095+2608:0+2608] <= intermediate[4095+2608:0+2608] + a; end
12'd2609: begin if(a[2609]==1) 
	 		intermediate[4095+2609:0+2609] <= intermediate[4095+2609:0+2609] + a; end
12'd2610: begin if(a[2610]==1) 
	 		intermediate[4095+2610:0+2610] <= intermediate[4095+2610:0+2610] + a; end
12'd2611: begin if(a[2611]==1) 
	 		intermediate[4095+2611:0+2611] <= intermediate[4095+2611:0+2611] + a; end
12'd2612: begin if(a[2612]==1) 
	 		intermediate[4095+2612:0+2612] <= intermediate[4095+2612:0+2612] + a; end
12'd2613: begin if(a[2613]==1) 
	 		intermediate[4095+2613:0+2613] <= intermediate[4095+2613:0+2613] + a; end
12'd2614: begin if(a[2614]==1) 
	 		intermediate[4095+2614:0+2614] <= intermediate[4095+2614:0+2614] + a; end
12'd2615: begin if(a[2615]==1) 
	 		intermediate[4095+2615:0+2615] <= intermediate[4095+2615:0+2615] + a; end
12'd2616: begin if(a[2616]==1) 
	 		intermediate[4095+2616:0+2616] <= intermediate[4095+2616:0+2616] + a; end
12'd2617: begin if(a[2617]==1) 
	 		intermediate[4095+2617:0+2617] <= intermediate[4095+2617:0+2617] + a; end
12'd2618: begin if(a[2618]==1) 
	 		intermediate[4095+2618:0+2618] <= intermediate[4095+2618:0+2618] + a; end
12'd2619: begin if(a[2619]==1) 
	 		intermediate[4095+2619:0+2619] <= intermediate[4095+2619:0+2619] + a; end
12'd2620: begin if(a[2620]==1) 
	 		intermediate[4095+2620:0+2620] <= intermediate[4095+2620:0+2620] + a; end
12'd2621: begin if(a[2621]==1) 
	 		intermediate[4095+2621:0+2621] <= intermediate[4095+2621:0+2621] + a; end
12'd2622: begin if(a[2622]==1) 
	 		intermediate[4095+2622:0+2622] <= intermediate[4095+2622:0+2622] + a; end
12'd2623: begin if(a[2623]==1) 
	 		intermediate[4095+2623:0+2623] <= intermediate[4095+2623:0+2623] + a; end
12'd2624: begin if(a[2624]==1) 
	 		intermediate[4095+2624:0+2624] <= intermediate[4095+2624:0+2624] + a; end
12'd2625: begin if(a[2625]==1) 
	 		intermediate[4095+2625:0+2625] <= intermediate[4095+2625:0+2625] + a; end
12'd2626: begin if(a[2626]==1) 
	 		intermediate[4095+2626:0+2626] <= intermediate[4095+2626:0+2626] + a; end
12'd2627: begin if(a[2627]==1) 
	 		intermediate[4095+2627:0+2627] <= intermediate[4095+2627:0+2627] + a; end
12'd2628: begin if(a[2628]==1) 
	 		intermediate[4095+2628:0+2628] <= intermediate[4095+2628:0+2628] + a; end
12'd2629: begin if(a[2629]==1) 
	 		intermediate[4095+2629:0+2629] <= intermediate[4095+2629:0+2629] + a; end
12'd2630: begin if(a[2630]==1) 
	 		intermediate[4095+2630:0+2630] <= intermediate[4095+2630:0+2630] + a; end
12'd2631: begin if(a[2631]==1) 
	 		intermediate[4095+2631:0+2631] <= intermediate[4095+2631:0+2631] + a; end
12'd2632: begin if(a[2632]==1) 
	 		intermediate[4095+2632:0+2632] <= intermediate[4095+2632:0+2632] + a; end
12'd2633: begin if(a[2633]==1) 
	 		intermediate[4095+2633:0+2633] <= intermediate[4095+2633:0+2633] + a; end
12'd2634: begin if(a[2634]==1) 
	 		intermediate[4095+2634:0+2634] <= intermediate[4095+2634:0+2634] + a; end
12'd2635: begin if(a[2635]==1) 
	 		intermediate[4095+2635:0+2635] <= intermediate[4095+2635:0+2635] + a; end
12'd2636: begin if(a[2636]==1) 
	 		intermediate[4095+2636:0+2636] <= intermediate[4095+2636:0+2636] + a; end
12'd2637: begin if(a[2637]==1) 
	 		intermediate[4095+2637:0+2637] <= intermediate[4095+2637:0+2637] + a; end
12'd2638: begin if(a[2638]==1) 
	 		intermediate[4095+2638:0+2638] <= intermediate[4095+2638:0+2638] + a; end
12'd2639: begin if(a[2639]==1) 
	 		intermediate[4095+2639:0+2639] <= intermediate[4095+2639:0+2639] + a; end
12'd2640: begin if(a[2640]==1) 
	 		intermediate[4095+2640:0+2640] <= intermediate[4095+2640:0+2640] + a; end
12'd2641: begin if(a[2641]==1) 
	 		intermediate[4095+2641:0+2641] <= intermediate[4095+2641:0+2641] + a; end
12'd2642: begin if(a[2642]==1) 
	 		intermediate[4095+2642:0+2642] <= intermediate[4095+2642:0+2642] + a; end
12'd2643: begin if(a[2643]==1) 
	 		intermediate[4095+2643:0+2643] <= intermediate[4095+2643:0+2643] + a; end
12'd2644: begin if(a[2644]==1) 
	 		intermediate[4095+2644:0+2644] <= intermediate[4095+2644:0+2644] + a; end
12'd2645: begin if(a[2645]==1) 
	 		intermediate[4095+2645:0+2645] <= intermediate[4095+2645:0+2645] + a; end
12'd2646: begin if(a[2646]==1) 
	 		intermediate[4095+2646:0+2646] <= intermediate[4095+2646:0+2646] + a; end
12'd2647: begin if(a[2647]==1) 
	 		intermediate[4095+2647:0+2647] <= intermediate[4095+2647:0+2647] + a; end
12'd2648: begin if(a[2648]==1) 
	 		intermediate[4095+2648:0+2648] <= intermediate[4095+2648:0+2648] + a; end
12'd2649: begin if(a[2649]==1) 
	 		intermediate[4095+2649:0+2649] <= intermediate[4095+2649:0+2649] + a; end
12'd2650: begin if(a[2650]==1) 
	 		intermediate[4095+2650:0+2650] <= intermediate[4095+2650:0+2650] + a; end
12'd2651: begin if(a[2651]==1) 
	 		intermediate[4095+2651:0+2651] <= intermediate[4095+2651:0+2651] + a; end
12'd2652: begin if(a[2652]==1) 
	 		intermediate[4095+2652:0+2652] <= intermediate[4095+2652:0+2652] + a; end
12'd2653: begin if(a[2653]==1) 
	 		intermediate[4095+2653:0+2653] <= intermediate[4095+2653:0+2653] + a; end
12'd2654: begin if(a[2654]==1) 
	 		intermediate[4095+2654:0+2654] <= intermediate[4095+2654:0+2654] + a; end
12'd2655: begin if(a[2655]==1) 
	 		intermediate[4095+2655:0+2655] <= intermediate[4095+2655:0+2655] + a; end
12'd2656: begin if(a[2656]==1) 
	 		intermediate[4095+2656:0+2656] <= intermediate[4095+2656:0+2656] + a; end
12'd2657: begin if(a[2657]==1) 
	 		intermediate[4095+2657:0+2657] <= intermediate[4095+2657:0+2657] + a; end
12'd2658: begin if(a[2658]==1) 
	 		intermediate[4095+2658:0+2658] <= intermediate[4095+2658:0+2658] + a; end
12'd2659: begin if(a[2659]==1) 
	 		intermediate[4095+2659:0+2659] <= intermediate[4095+2659:0+2659] + a; end
12'd2660: begin if(a[2660]==1) 
	 		intermediate[4095+2660:0+2660] <= intermediate[4095+2660:0+2660] + a; end
12'd2661: begin if(a[2661]==1) 
	 		intermediate[4095+2661:0+2661] <= intermediate[4095+2661:0+2661] + a; end
12'd2662: begin if(a[2662]==1) 
	 		intermediate[4095+2662:0+2662] <= intermediate[4095+2662:0+2662] + a; end
12'd2663: begin if(a[2663]==1) 
	 		intermediate[4095+2663:0+2663] <= intermediate[4095+2663:0+2663] + a; end
12'd2664: begin if(a[2664]==1) 
	 		intermediate[4095+2664:0+2664] <= intermediate[4095+2664:0+2664] + a; end
12'd2665: begin if(a[2665]==1) 
	 		intermediate[4095+2665:0+2665] <= intermediate[4095+2665:0+2665] + a; end
12'd2666: begin if(a[2666]==1) 
	 		intermediate[4095+2666:0+2666] <= intermediate[4095+2666:0+2666] + a; end
12'd2667: begin if(a[2667]==1) 
	 		intermediate[4095+2667:0+2667] <= intermediate[4095+2667:0+2667] + a; end
12'd2668: begin if(a[2668]==1) 
	 		intermediate[4095+2668:0+2668] <= intermediate[4095+2668:0+2668] + a; end
12'd2669: begin if(a[2669]==1) 
	 		intermediate[4095+2669:0+2669] <= intermediate[4095+2669:0+2669] + a; end
12'd2670: begin if(a[2670]==1) 
	 		intermediate[4095+2670:0+2670] <= intermediate[4095+2670:0+2670] + a; end
12'd2671: begin if(a[2671]==1) 
	 		intermediate[4095+2671:0+2671] <= intermediate[4095+2671:0+2671] + a; end
12'd2672: begin if(a[2672]==1) 
	 		intermediate[4095+2672:0+2672] <= intermediate[4095+2672:0+2672] + a; end
12'd2673: begin if(a[2673]==1) 
	 		intermediate[4095+2673:0+2673] <= intermediate[4095+2673:0+2673] + a; end
12'd2674: begin if(a[2674]==1) 
	 		intermediate[4095+2674:0+2674] <= intermediate[4095+2674:0+2674] + a; end
12'd2675: begin if(a[2675]==1) 
	 		intermediate[4095+2675:0+2675] <= intermediate[4095+2675:0+2675] + a; end
12'd2676: begin if(a[2676]==1) 
	 		intermediate[4095+2676:0+2676] <= intermediate[4095+2676:0+2676] + a; end
12'd2677: begin if(a[2677]==1) 
	 		intermediate[4095+2677:0+2677] <= intermediate[4095+2677:0+2677] + a; end
12'd2678: begin if(a[2678]==1) 
	 		intermediate[4095+2678:0+2678] <= intermediate[4095+2678:0+2678] + a; end
12'd2679: begin if(a[2679]==1) 
	 		intermediate[4095+2679:0+2679] <= intermediate[4095+2679:0+2679] + a; end
12'd2680: begin if(a[2680]==1) 
	 		intermediate[4095+2680:0+2680] <= intermediate[4095+2680:0+2680] + a; end
12'd2681: begin if(a[2681]==1) 
	 		intermediate[4095+2681:0+2681] <= intermediate[4095+2681:0+2681] + a; end
12'd2682: begin if(a[2682]==1) 
	 		intermediate[4095+2682:0+2682] <= intermediate[4095+2682:0+2682] + a; end
12'd2683: begin if(a[2683]==1) 
	 		intermediate[4095+2683:0+2683] <= intermediate[4095+2683:0+2683] + a; end
12'd2684: begin if(a[2684]==1) 
	 		intermediate[4095+2684:0+2684] <= intermediate[4095+2684:0+2684] + a; end
12'd2685: begin if(a[2685]==1) 
	 		intermediate[4095+2685:0+2685] <= intermediate[4095+2685:0+2685] + a; end
12'd2686: begin if(a[2686]==1) 
	 		intermediate[4095+2686:0+2686] <= intermediate[4095+2686:0+2686] + a; end
12'd2687: begin if(a[2687]==1) 
	 		intermediate[4095+2687:0+2687] <= intermediate[4095+2687:0+2687] + a; end
12'd2688: begin if(a[2688]==1) 
	 		intermediate[4095+2688:0+2688] <= intermediate[4095+2688:0+2688] + a; end
12'd2689: begin if(a[2689]==1) 
	 		intermediate[4095+2689:0+2689] <= intermediate[4095+2689:0+2689] + a; end
12'd2690: begin if(a[2690]==1) 
	 		intermediate[4095+2690:0+2690] <= intermediate[4095+2690:0+2690] + a; end
12'd2691: begin if(a[2691]==1) 
	 		intermediate[4095+2691:0+2691] <= intermediate[4095+2691:0+2691] + a; end
12'd2692: begin if(a[2692]==1) 
	 		intermediate[4095+2692:0+2692] <= intermediate[4095+2692:0+2692] + a; end
12'd2693: begin if(a[2693]==1) 
	 		intermediate[4095+2693:0+2693] <= intermediate[4095+2693:0+2693] + a; end
12'd2694: begin if(a[2694]==1) 
	 		intermediate[4095+2694:0+2694] <= intermediate[4095+2694:0+2694] + a; end
12'd2695: begin if(a[2695]==1) 
	 		intermediate[4095+2695:0+2695] <= intermediate[4095+2695:0+2695] + a; end
12'd2696: begin if(a[2696]==1) 
	 		intermediate[4095+2696:0+2696] <= intermediate[4095+2696:0+2696] + a; end
12'd2697: begin if(a[2697]==1) 
	 		intermediate[4095+2697:0+2697] <= intermediate[4095+2697:0+2697] + a; end
12'd2698: begin if(a[2698]==1) 
	 		intermediate[4095+2698:0+2698] <= intermediate[4095+2698:0+2698] + a; end
12'd2699: begin if(a[2699]==1) 
	 		intermediate[4095+2699:0+2699] <= intermediate[4095+2699:0+2699] + a; end
12'd2700: begin if(a[2700]==1) 
	 		intermediate[4095+2700:0+2700] <= intermediate[4095+2700:0+2700] + a; end
12'd2701: begin if(a[2701]==1) 
	 		intermediate[4095+2701:0+2701] <= intermediate[4095+2701:0+2701] + a; end
12'd2702: begin if(a[2702]==1) 
	 		intermediate[4095+2702:0+2702] <= intermediate[4095+2702:0+2702] + a; end
12'd2703: begin if(a[2703]==1) 
	 		intermediate[4095+2703:0+2703] <= intermediate[4095+2703:0+2703] + a; end
12'd2704: begin if(a[2704]==1) 
	 		intermediate[4095+2704:0+2704] <= intermediate[4095+2704:0+2704] + a; end
12'd2705: begin if(a[2705]==1) 
	 		intermediate[4095+2705:0+2705] <= intermediate[4095+2705:0+2705] + a; end
12'd2706: begin if(a[2706]==1) 
	 		intermediate[4095+2706:0+2706] <= intermediate[4095+2706:0+2706] + a; end
12'd2707: begin if(a[2707]==1) 
	 		intermediate[4095+2707:0+2707] <= intermediate[4095+2707:0+2707] + a; end
12'd2708: begin if(a[2708]==1) 
	 		intermediate[4095+2708:0+2708] <= intermediate[4095+2708:0+2708] + a; end
12'd2709: begin if(a[2709]==1) 
	 		intermediate[4095+2709:0+2709] <= intermediate[4095+2709:0+2709] + a; end
12'd2710: begin if(a[2710]==1) 
	 		intermediate[4095+2710:0+2710] <= intermediate[4095+2710:0+2710] + a; end
12'd2711: begin if(a[2711]==1) 
	 		intermediate[4095+2711:0+2711] <= intermediate[4095+2711:0+2711] + a; end
12'd2712: begin if(a[2712]==1) 
	 		intermediate[4095+2712:0+2712] <= intermediate[4095+2712:0+2712] + a; end
12'd2713: begin if(a[2713]==1) 
	 		intermediate[4095+2713:0+2713] <= intermediate[4095+2713:0+2713] + a; end
12'd2714: begin if(a[2714]==1) 
	 		intermediate[4095+2714:0+2714] <= intermediate[4095+2714:0+2714] + a; end
12'd2715: begin if(a[2715]==1) 
	 		intermediate[4095+2715:0+2715] <= intermediate[4095+2715:0+2715] + a; end
12'd2716: begin if(a[2716]==1) 
	 		intermediate[4095+2716:0+2716] <= intermediate[4095+2716:0+2716] + a; end
12'd2717: begin if(a[2717]==1) 
	 		intermediate[4095+2717:0+2717] <= intermediate[4095+2717:0+2717] + a; end
12'd2718: begin if(a[2718]==1) 
	 		intermediate[4095+2718:0+2718] <= intermediate[4095+2718:0+2718] + a; end
12'd2719: begin if(a[2719]==1) 
	 		intermediate[4095+2719:0+2719] <= intermediate[4095+2719:0+2719] + a; end
12'd2720: begin if(a[2720]==1) 
	 		intermediate[4095+2720:0+2720] <= intermediate[4095+2720:0+2720] + a; end
12'd2721: begin if(a[2721]==1) 
	 		intermediate[4095+2721:0+2721] <= intermediate[4095+2721:0+2721] + a; end
12'd2722: begin if(a[2722]==1) 
	 		intermediate[4095+2722:0+2722] <= intermediate[4095+2722:0+2722] + a; end
12'd2723: begin if(a[2723]==1) 
	 		intermediate[4095+2723:0+2723] <= intermediate[4095+2723:0+2723] + a; end
12'd2724: begin if(a[2724]==1) 
	 		intermediate[4095+2724:0+2724] <= intermediate[4095+2724:0+2724] + a; end
12'd2725: begin if(a[2725]==1) 
	 		intermediate[4095+2725:0+2725] <= intermediate[4095+2725:0+2725] + a; end
12'd2726: begin if(a[2726]==1) 
	 		intermediate[4095+2726:0+2726] <= intermediate[4095+2726:0+2726] + a; end
12'd2727: begin if(a[2727]==1) 
	 		intermediate[4095+2727:0+2727] <= intermediate[4095+2727:0+2727] + a; end
12'd2728: begin if(a[2728]==1) 
	 		intermediate[4095+2728:0+2728] <= intermediate[4095+2728:0+2728] + a; end
12'd2729: begin if(a[2729]==1) 
	 		intermediate[4095+2729:0+2729] <= intermediate[4095+2729:0+2729] + a; end
12'd2730: begin if(a[2730]==1) 
	 		intermediate[4095+2730:0+2730] <= intermediate[4095+2730:0+2730] + a; end
12'd2731: begin if(a[2731]==1) 
	 		intermediate[4095+2731:0+2731] <= intermediate[4095+2731:0+2731] + a; end
12'd2732: begin if(a[2732]==1) 
	 		intermediate[4095+2732:0+2732] <= intermediate[4095+2732:0+2732] + a; end
12'd2733: begin if(a[2733]==1) 
	 		intermediate[4095+2733:0+2733] <= intermediate[4095+2733:0+2733] + a; end
12'd2734: begin if(a[2734]==1) 
	 		intermediate[4095+2734:0+2734] <= intermediate[4095+2734:0+2734] + a; end
12'd2735: begin if(a[2735]==1) 
	 		intermediate[4095+2735:0+2735] <= intermediate[4095+2735:0+2735] + a; end
12'd2736: begin if(a[2736]==1) 
	 		intermediate[4095+2736:0+2736] <= intermediate[4095+2736:0+2736] + a; end
12'd2737: begin if(a[2737]==1) 
	 		intermediate[4095+2737:0+2737] <= intermediate[4095+2737:0+2737] + a; end
12'd2738: begin if(a[2738]==1) 
	 		intermediate[4095+2738:0+2738] <= intermediate[4095+2738:0+2738] + a; end
12'd2739: begin if(a[2739]==1) 
	 		intermediate[4095+2739:0+2739] <= intermediate[4095+2739:0+2739] + a; end
12'd2740: begin if(a[2740]==1) 
	 		intermediate[4095+2740:0+2740] <= intermediate[4095+2740:0+2740] + a; end
12'd2741: begin if(a[2741]==1) 
	 		intermediate[4095+2741:0+2741] <= intermediate[4095+2741:0+2741] + a; end
12'd2742: begin if(a[2742]==1) 
	 		intermediate[4095+2742:0+2742] <= intermediate[4095+2742:0+2742] + a; end
12'd2743: begin if(a[2743]==1) 
	 		intermediate[4095+2743:0+2743] <= intermediate[4095+2743:0+2743] + a; end
12'd2744: begin if(a[2744]==1) 
	 		intermediate[4095+2744:0+2744] <= intermediate[4095+2744:0+2744] + a; end
12'd2745: begin if(a[2745]==1) 
	 		intermediate[4095+2745:0+2745] <= intermediate[4095+2745:0+2745] + a; end
12'd2746: begin if(a[2746]==1) 
	 		intermediate[4095+2746:0+2746] <= intermediate[4095+2746:0+2746] + a; end
12'd2747: begin if(a[2747]==1) 
	 		intermediate[4095+2747:0+2747] <= intermediate[4095+2747:0+2747] + a; end
12'd2748: begin if(a[2748]==1) 
	 		intermediate[4095+2748:0+2748] <= intermediate[4095+2748:0+2748] + a; end
12'd2749: begin if(a[2749]==1) 
	 		intermediate[4095+2749:0+2749] <= intermediate[4095+2749:0+2749] + a; end
12'd2750: begin if(a[2750]==1) 
	 		intermediate[4095+2750:0+2750] <= intermediate[4095+2750:0+2750] + a; end
12'd2751: begin if(a[2751]==1) 
	 		intermediate[4095+2751:0+2751] <= intermediate[4095+2751:0+2751] + a; end
12'd2752: begin if(a[2752]==1) 
	 		intermediate[4095+2752:0+2752] <= intermediate[4095+2752:0+2752] + a; end
12'd2753: begin if(a[2753]==1) 
	 		intermediate[4095+2753:0+2753] <= intermediate[4095+2753:0+2753] + a; end
12'd2754: begin if(a[2754]==1) 
	 		intermediate[4095+2754:0+2754] <= intermediate[4095+2754:0+2754] + a; end
12'd2755: begin if(a[2755]==1) 
	 		intermediate[4095+2755:0+2755] <= intermediate[4095+2755:0+2755] + a; end
12'd2756: begin if(a[2756]==1) 
	 		intermediate[4095+2756:0+2756] <= intermediate[4095+2756:0+2756] + a; end
12'd2757: begin if(a[2757]==1) 
	 		intermediate[4095+2757:0+2757] <= intermediate[4095+2757:0+2757] + a; end
12'd2758: begin if(a[2758]==1) 
	 		intermediate[4095+2758:0+2758] <= intermediate[4095+2758:0+2758] + a; end
12'd2759: begin if(a[2759]==1) 
	 		intermediate[4095+2759:0+2759] <= intermediate[4095+2759:0+2759] + a; end
12'd2760: begin if(a[2760]==1) 
	 		intermediate[4095+2760:0+2760] <= intermediate[4095+2760:0+2760] + a; end
12'd2761: begin if(a[2761]==1) 
	 		intermediate[4095+2761:0+2761] <= intermediate[4095+2761:0+2761] + a; end
12'd2762: begin if(a[2762]==1) 
	 		intermediate[4095+2762:0+2762] <= intermediate[4095+2762:0+2762] + a; end
12'd2763: begin if(a[2763]==1) 
	 		intermediate[4095+2763:0+2763] <= intermediate[4095+2763:0+2763] + a; end
12'd2764: begin if(a[2764]==1) 
	 		intermediate[4095+2764:0+2764] <= intermediate[4095+2764:0+2764] + a; end
12'd2765: begin if(a[2765]==1) 
	 		intermediate[4095+2765:0+2765] <= intermediate[4095+2765:0+2765] + a; end
12'd2766: begin if(a[2766]==1) 
	 		intermediate[4095+2766:0+2766] <= intermediate[4095+2766:0+2766] + a; end
12'd2767: begin if(a[2767]==1) 
	 		intermediate[4095+2767:0+2767] <= intermediate[4095+2767:0+2767] + a; end
12'd2768: begin if(a[2768]==1) 
	 		intermediate[4095+2768:0+2768] <= intermediate[4095+2768:0+2768] + a; end
12'd2769: begin if(a[2769]==1) 
	 		intermediate[4095+2769:0+2769] <= intermediate[4095+2769:0+2769] + a; end
12'd2770: begin if(a[2770]==1) 
	 		intermediate[4095+2770:0+2770] <= intermediate[4095+2770:0+2770] + a; end
12'd2771: begin if(a[2771]==1) 
	 		intermediate[4095+2771:0+2771] <= intermediate[4095+2771:0+2771] + a; end
12'd2772: begin if(a[2772]==1) 
	 		intermediate[4095+2772:0+2772] <= intermediate[4095+2772:0+2772] + a; end
12'd2773: begin if(a[2773]==1) 
	 		intermediate[4095+2773:0+2773] <= intermediate[4095+2773:0+2773] + a; end
12'd2774: begin if(a[2774]==1) 
	 		intermediate[4095+2774:0+2774] <= intermediate[4095+2774:0+2774] + a; end
12'd2775: begin if(a[2775]==1) 
	 		intermediate[4095+2775:0+2775] <= intermediate[4095+2775:0+2775] + a; end
12'd2776: begin if(a[2776]==1) 
	 		intermediate[4095+2776:0+2776] <= intermediate[4095+2776:0+2776] + a; end
12'd2777: begin if(a[2777]==1) 
	 		intermediate[4095+2777:0+2777] <= intermediate[4095+2777:0+2777] + a; end
12'd2778: begin if(a[2778]==1) 
	 		intermediate[4095+2778:0+2778] <= intermediate[4095+2778:0+2778] + a; end
12'd2779: begin if(a[2779]==1) 
	 		intermediate[4095+2779:0+2779] <= intermediate[4095+2779:0+2779] + a; end
12'd2780: begin if(a[2780]==1) 
	 		intermediate[4095+2780:0+2780] <= intermediate[4095+2780:0+2780] + a; end
12'd2781: begin if(a[2781]==1) 
	 		intermediate[4095+2781:0+2781] <= intermediate[4095+2781:0+2781] + a; end
12'd2782: begin if(a[2782]==1) 
	 		intermediate[4095+2782:0+2782] <= intermediate[4095+2782:0+2782] + a; end
12'd2783: begin if(a[2783]==1) 
	 		intermediate[4095+2783:0+2783] <= intermediate[4095+2783:0+2783] + a; end
12'd2784: begin if(a[2784]==1) 
	 		intermediate[4095+2784:0+2784] <= intermediate[4095+2784:0+2784] + a; end
12'd2785: begin if(a[2785]==1) 
	 		intermediate[4095+2785:0+2785] <= intermediate[4095+2785:0+2785] + a; end
12'd2786: begin if(a[2786]==1) 
	 		intermediate[4095+2786:0+2786] <= intermediate[4095+2786:0+2786] + a; end
12'd2787: begin if(a[2787]==1) 
	 		intermediate[4095+2787:0+2787] <= intermediate[4095+2787:0+2787] + a; end
12'd2788: begin if(a[2788]==1) 
	 		intermediate[4095+2788:0+2788] <= intermediate[4095+2788:0+2788] + a; end
12'd2789: begin if(a[2789]==1) 
	 		intermediate[4095+2789:0+2789] <= intermediate[4095+2789:0+2789] + a; end
12'd2790: begin if(a[2790]==1) 
	 		intermediate[4095+2790:0+2790] <= intermediate[4095+2790:0+2790] + a; end
12'd2791: begin if(a[2791]==1) 
	 		intermediate[4095+2791:0+2791] <= intermediate[4095+2791:0+2791] + a; end
12'd2792: begin if(a[2792]==1) 
	 		intermediate[4095+2792:0+2792] <= intermediate[4095+2792:0+2792] + a; end
12'd2793: begin if(a[2793]==1) 
	 		intermediate[4095+2793:0+2793] <= intermediate[4095+2793:0+2793] + a; end
12'd2794: begin if(a[2794]==1) 
	 		intermediate[4095+2794:0+2794] <= intermediate[4095+2794:0+2794] + a; end
12'd2795: begin if(a[2795]==1) 
	 		intermediate[4095+2795:0+2795] <= intermediate[4095+2795:0+2795] + a; end
12'd2796: begin if(a[2796]==1) 
	 		intermediate[4095+2796:0+2796] <= intermediate[4095+2796:0+2796] + a; end
12'd2797: begin if(a[2797]==1) 
	 		intermediate[4095+2797:0+2797] <= intermediate[4095+2797:0+2797] + a; end
12'd2798: begin if(a[2798]==1) 
	 		intermediate[4095+2798:0+2798] <= intermediate[4095+2798:0+2798] + a; end
12'd2799: begin if(a[2799]==1) 
	 		intermediate[4095+2799:0+2799] <= intermediate[4095+2799:0+2799] + a; end
12'd2800: begin if(a[2800]==1) 
	 		intermediate[4095+2800:0+2800] <= intermediate[4095+2800:0+2800] + a; end
12'd2801: begin if(a[2801]==1) 
	 		intermediate[4095+2801:0+2801] <= intermediate[4095+2801:0+2801] + a; end
12'd2802: begin if(a[2802]==1) 
	 		intermediate[4095+2802:0+2802] <= intermediate[4095+2802:0+2802] + a; end
12'd2803: begin if(a[2803]==1) 
	 		intermediate[4095+2803:0+2803] <= intermediate[4095+2803:0+2803] + a; end
12'd2804: begin if(a[2804]==1) 
	 		intermediate[4095+2804:0+2804] <= intermediate[4095+2804:0+2804] + a; end
12'd2805: begin if(a[2805]==1) 
	 		intermediate[4095+2805:0+2805] <= intermediate[4095+2805:0+2805] + a; end
12'd2806: begin if(a[2806]==1) 
	 		intermediate[4095+2806:0+2806] <= intermediate[4095+2806:0+2806] + a; end
12'd2807: begin if(a[2807]==1) 
	 		intermediate[4095+2807:0+2807] <= intermediate[4095+2807:0+2807] + a; end
12'd2808: begin if(a[2808]==1) 
	 		intermediate[4095+2808:0+2808] <= intermediate[4095+2808:0+2808] + a; end
12'd2809: begin if(a[2809]==1) 
	 		intermediate[4095+2809:0+2809] <= intermediate[4095+2809:0+2809] + a; end
12'd2810: begin if(a[2810]==1) 
	 		intermediate[4095+2810:0+2810] <= intermediate[4095+2810:0+2810] + a; end
12'd2811: begin if(a[2811]==1) 
	 		intermediate[4095+2811:0+2811] <= intermediate[4095+2811:0+2811] + a; end
12'd2812: begin if(a[2812]==1) 
	 		intermediate[4095+2812:0+2812] <= intermediate[4095+2812:0+2812] + a; end
12'd2813: begin if(a[2813]==1) 
	 		intermediate[4095+2813:0+2813] <= intermediate[4095+2813:0+2813] + a; end
12'd2814: begin if(a[2814]==1) 
	 		intermediate[4095+2814:0+2814] <= intermediate[4095+2814:0+2814] + a; end
12'd2815: begin if(a[2815]==1) 
	 		intermediate[4095+2815:0+2815] <= intermediate[4095+2815:0+2815] + a; end
12'd2816: begin if(a[2816]==1) 
	 		intermediate[4095+2816:0+2816] <= intermediate[4095+2816:0+2816] + a; end
12'd2817: begin if(a[2817]==1) 
	 		intermediate[4095+2817:0+2817] <= intermediate[4095+2817:0+2817] + a; end
12'd2818: begin if(a[2818]==1) 
	 		intermediate[4095+2818:0+2818] <= intermediate[4095+2818:0+2818] + a; end
12'd2819: begin if(a[2819]==1) 
	 		intermediate[4095+2819:0+2819] <= intermediate[4095+2819:0+2819] + a; end
12'd2820: begin if(a[2820]==1) 
	 		intermediate[4095+2820:0+2820] <= intermediate[4095+2820:0+2820] + a; end
12'd2821: begin if(a[2821]==1) 
	 		intermediate[4095+2821:0+2821] <= intermediate[4095+2821:0+2821] + a; end
12'd2822: begin if(a[2822]==1) 
	 		intermediate[4095+2822:0+2822] <= intermediate[4095+2822:0+2822] + a; end
12'd2823: begin if(a[2823]==1) 
	 		intermediate[4095+2823:0+2823] <= intermediate[4095+2823:0+2823] + a; end
12'd2824: begin if(a[2824]==1) 
	 		intermediate[4095+2824:0+2824] <= intermediate[4095+2824:0+2824] + a; end
12'd2825: begin if(a[2825]==1) 
	 		intermediate[4095+2825:0+2825] <= intermediate[4095+2825:0+2825] + a; end
12'd2826: begin if(a[2826]==1) 
	 		intermediate[4095+2826:0+2826] <= intermediate[4095+2826:0+2826] + a; end
12'd2827: begin if(a[2827]==1) 
	 		intermediate[4095+2827:0+2827] <= intermediate[4095+2827:0+2827] + a; end
12'd2828: begin if(a[2828]==1) 
	 		intermediate[4095+2828:0+2828] <= intermediate[4095+2828:0+2828] + a; end
12'd2829: begin if(a[2829]==1) 
	 		intermediate[4095+2829:0+2829] <= intermediate[4095+2829:0+2829] + a; end
12'd2830: begin if(a[2830]==1) 
	 		intermediate[4095+2830:0+2830] <= intermediate[4095+2830:0+2830] + a; end
12'd2831: begin if(a[2831]==1) 
	 		intermediate[4095+2831:0+2831] <= intermediate[4095+2831:0+2831] + a; end
12'd2832: begin if(a[2832]==1) 
	 		intermediate[4095+2832:0+2832] <= intermediate[4095+2832:0+2832] + a; end
12'd2833: begin if(a[2833]==1) 
	 		intermediate[4095+2833:0+2833] <= intermediate[4095+2833:0+2833] + a; end
12'd2834: begin if(a[2834]==1) 
	 		intermediate[4095+2834:0+2834] <= intermediate[4095+2834:0+2834] + a; end
12'd2835: begin if(a[2835]==1) 
	 		intermediate[4095+2835:0+2835] <= intermediate[4095+2835:0+2835] + a; end
12'd2836: begin if(a[2836]==1) 
	 		intermediate[4095+2836:0+2836] <= intermediate[4095+2836:0+2836] + a; end
12'd2837: begin if(a[2837]==1) 
	 		intermediate[4095+2837:0+2837] <= intermediate[4095+2837:0+2837] + a; end
12'd2838: begin if(a[2838]==1) 
	 		intermediate[4095+2838:0+2838] <= intermediate[4095+2838:0+2838] + a; end
12'd2839: begin if(a[2839]==1) 
	 		intermediate[4095+2839:0+2839] <= intermediate[4095+2839:0+2839] + a; end
12'd2840: begin if(a[2840]==1) 
	 		intermediate[4095+2840:0+2840] <= intermediate[4095+2840:0+2840] + a; end
12'd2841: begin if(a[2841]==1) 
	 		intermediate[4095+2841:0+2841] <= intermediate[4095+2841:0+2841] + a; end
12'd2842: begin if(a[2842]==1) 
	 		intermediate[4095+2842:0+2842] <= intermediate[4095+2842:0+2842] + a; end
12'd2843: begin if(a[2843]==1) 
	 		intermediate[4095+2843:0+2843] <= intermediate[4095+2843:0+2843] + a; end
12'd2844: begin if(a[2844]==1) 
	 		intermediate[4095+2844:0+2844] <= intermediate[4095+2844:0+2844] + a; end
12'd2845: begin if(a[2845]==1) 
	 		intermediate[4095+2845:0+2845] <= intermediate[4095+2845:0+2845] + a; end
12'd2846: begin if(a[2846]==1) 
	 		intermediate[4095+2846:0+2846] <= intermediate[4095+2846:0+2846] + a; end
12'd2847: begin if(a[2847]==1) 
	 		intermediate[4095+2847:0+2847] <= intermediate[4095+2847:0+2847] + a; end
12'd2848: begin if(a[2848]==1) 
	 		intermediate[4095+2848:0+2848] <= intermediate[4095+2848:0+2848] + a; end
12'd2849: begin if(a[2849]==1) 
	 		intermediate[4095+2849:0+2849] <= intermediate[4095+2849:0+2849] + a; end
12'd2850: begin if(a[2850]==1) 
	 		intermediate[4095+2850:0+2850] <= intermediate[4095+2850:0+2850] + a; end
12'd2851: begin if(a[2851]==1) 
	 		intermediate[4095+2851:0+2851] <= intermediate[4095+2851:0+2851] + a; end
12'd2852: begin if(a[2852]==1) 
	 		intermediate[4095+2852:0+2852] <= intermediate[4095+2852:0+2852] + a; end
12'd2853: begin if(a[2853]==1) 
	 		intermediate[4095+2853:0+2853] <= intermediate[4095+2853:0+2853] + a; end
12'd2854: begin if(a[2854]==1) 
	 		intermediate[4095+2854:0+2854] <= intermediate[4095+2854:0+2854] + a; end
12'd2855: begin if(a[2855]==1) 
	 		intermediate[4095+2855:0+2855] <= intermediate[4095+2855:0+2855] + a; end
12'd2856: begin if(a[2856]==1) 
	 		intermediate[4095+2856:0+2856] <= intermediate[4095+2856:0+2856] + a; end
12'd2857: begin if(a[2857]==1) 
	 		intermediate[4095+2857:0+2857] <= intermediate[4095+2857:0+2857] + a; end
12'd2858: begin if(a[2858]==1) 
	 		intermediate[4095+2858:0+2858] <= intermediate[4095+2858:0+2858] + a; end
12'd2859: begin if(a[2859]==1) 
	 		intermediate[4095+2859:0+2859] <= intermediate[4095+2859:0+2859] + a; end
12'd2860: begin if(a[2860]==1) 
	 		intermediate[4095+2860:0+2860] <= intermediate[4095+2860:0+2860] + a; end
12'd2861: begin if(a[2861]==1) 
	 		intermediate[4095+2861:0+2861] <= intermediate[4095+2861:0+2861] + a; end
12'd2862: begin if(a[2862]==1) 
	 		intermediate[4095+2862:0+2862] <= intermediate[4095+2862:0+2862] + a; end
12'd2863: begin if(a[2863]==1) 
	 		intermediate[4095+2863:0+2863] <= intermediate[4095+2863:0+2863] + a; end
12'd2864: begin if(a[2864]==1) 
	 		intermediate[4095+2864:0+2864] <= intermediate[4095+2864:0+2864] + a; end
12'd2865: begin if(a[2865]==1) 
	 		intermediate[4095+2865:0+2865] <= intermediate[4095+2865:0+2865] + a; end
12'd2866: begin if(a[2866]==1) 
	 		intermediate[4095+2866:0+2866] <= intermediate[4095+2866:0+2866] + a; end
12'd2867: begin if(a[2867]==1) 
	 		intermediate[4095+2867:0+2867] <= intermediate[4095+2867:0+2867] + a; end
12'd2868: begin if(a[2868]==1) 
	 		intermediate[4095+2868:0+2868] <= intermediate[4095+2868:0+2868] + a; end
12'd2869: begin if(a[2869]==1) 
	 		intermediate[4095+2869:0+2869] <= intermediate[4095+2869:0+2869] + a; end
12'd2870: begin if(a[2870]==1) 
	 		intermediate[4095+2870:0+2870] <= intermediate[4095+2870:0+2870] + a; end
12'd2871: begin if(a[2871]==1) 
	 		intermediate[4095+2871:0+2871] <= intermediate[4095+2871:0+2871] + a; end
12'd2872: begin if(a[2872]==1) 
	 		intermediate[4095+2872:0+2872] <= intermediate[4095+2872:0+2872] + a; end
12'd2873: begin if(a[2873]==1) 
	 		intermediate[4095+2873:0+2873] <= intermediate[4095+2873:0+2873] + a; end
12'd2874: begin if(a[2874]==1) 
	 		intermediate[4095+2874:0+2874] <= intermediate[4095+2874:0+2874] + a; end
12'd2875: begin if(a[2875]==1) 
	 		intermediate[4095+2875:0+2875] <= intermediate[4095+2875:0+2875] + a; end
12'd2876: begin if(a[2876]==1) 
	 		intermediate[4095+2876:0+2876] <= intermediate[4095+2876:0+2876] + a; end
12'd2877: begin if(a[2877]==1) 
	 		intermediate[4095+2877:0+2877] <= intermediate[4095+2877:0+2877] + a; end
12'd2878: begin if(a[2878]==1) 
	 		intermediate[4095+2878:0+2878] <= intermediate[4095+2878:0+2878] + a; end
12'd2879: begin if(a[2879]==1) 
	 		intermediate[4095+2879:0+2879] <= intermediate[4095+2879:0+2879] + a; end
12'd2880: begin if(a[2880]==1) 
	 		intermediate[4095+2880:0+2880] <= intermediate[4095+2880:0+2880] + a; end
12'd2881: begin if(a[2881]==1) 
	 		intermediate[4095+2881:0+2881] <= intermediate[4095+2881:0+2881] + a; end
12'd2882: begin if(a[2882]==1) 
	 		intermediate[4095+2882:0+2882] <= intermediate[4095+2882:0+2882] + a; end
12'd2883: begin if(a[2883]==1) 
	 		intermediate[4095+2883:0+2883] <= intermediate[4095+2883:0+2883] + a; end
12'd2884: begin if(a[2884]==1) 
	 		intermediate[4095+2884:0+2884] <= intermediate[4095+2884:0+2884] + a; end
12'd2885: begin if(a[2885]==1) 
	 		intermediate[4095+2885:0+2885] <= intermediate[4095+2885:0+2885] + a; end
12'd2886: begin if(a[2886]==1) 
	 		intermediate[4095+2886:0+2886] <= intermediate[4095+2886:0+2886] + a; end
12'd2887: begin if(a[2887]==1) 
	 		intermediate[4095+2887:0+2887] <= intermediate[4095+2887:0+2887] + a; end
12'd2888: begin if(a[2888]==1) 
	 		intermediate[4095+2888:0+2888] <= intermediate[4095+2888:0+2888] + a; end
12'd2889: begin if(a[2889]==1) 
	 		intermediate[4095+2889:0+2889] <= intermediate[4095+2889:0+2889] + a; end
12'd2890: begin if(a[2890]==1) 
	 		intermediate[4095+2890:0+2890] <= intermediate[4095+2890:0+2890] + a; end
12'd2891: begin if(a[2891]==1) 
	 		intermediate[4095+2891:0+2891] <= intermediate[4095+2891:0+2891] + a; end
12'd2892: begin if(a[2892]==1) 
	 		intermediate[4095+2892:0+2892] <= intermediate[4095+2892:0+2892] + a; end
12'd2893: begin if(a[2893]==1) 
	 		intermediate[4095+2893:0+2893] <= intermediate[4095+2893:0+2893] + a; end
12'd2894: begin if(a[2894]==1) 
	 		intermediate[4095+2894:0+2894] <= intermediate[4095+2894:0+2894] + a; end
12'd2895: begin if(a[2895]==1) 
	 		intermediate[4095+2895:0+2895] <= intermediate[4095+2895:0+2895] + a; end
12'd2896: begin if(a[2896]==1) 
	 		intermediate[4095+2896:0+2896] <= intermediate[4095+2896:0+2896] + a; end
12'd2897: begin if(a[2897]==1) 
	 		intermediate[4095+2897:0+2897] <= intermediate[4095+2897:0+2897] + a; end
12'd2898: begin if(a[2898]==1) 
	 		intermediate[4095+2898:0+2898] <= intermediate[4095+2898:0+2898] + a; end
12'd2899: begin if(a[2899]==1) 
	 		intermediate[4095+2899:0+2899] <= intermediate[4095+2899:0+2899] + a; end
12'd2900: begin if(a[2900]==1) 
	 		intermediate[4095+2900:0+2900] <= intermediate[4095+2900:0+2900] + a; end
12'd2901: begin if(a[2901]==1) 
	 		intermediate[4095+2901:0+2901] <= intermediate[4095+2901:0+2901] + a; end
12'd2902: begin if(a[2902]==1) 
	 		intermediate[4095+2902:0+2902] <= intermediate[4095+2902:0+2902] + a; end
12'd2903: begin if(a[2903]==1) 
	 		intermediate[4095+2903:0+2903] <= intermediate[4095+2903:0+2903] + a; end
12'd2904: begin if(a[2904]==1) 
	 		intermediate[4095+2904:0+2904] <= intermediate[4095+2904:0+2904] + a; end
12'd2905: begin if(a[2905]==1) 
	 		intermediate[4095+2905:0+2905] <= intermediate[4095+2905:0+2905] + a; end
12'd2906: begin if(a[2906]==1) 
	 		intermediate[4095+2906:0+2906] <= intermediate[4095+2906:0+2906] + a; end
12'd2907: begin if(a[2907]==1) 
	 		intermediate[4095+2907:0+2907] <= intermediate[4095+2907:0+2907] + a; end
12'd2908: begin if(a[2908]==1) 
	 		intermediate[4095+2908:0+2908] <= intermediate[4095+2908:0+2908] + a; end
12'd2909: begin if(a[2909]==1) 
	 		intermediate[4095+2909:0+2909] <= intermediate[4095+2909:0+2909] + a; end
12'd2910: begin if(a[2910]==1) 
	 		intermediate[4095+2910:0+2910] <= intermediate[4095+2910:0+2910] + a; end
12'd2911: begin if(a[2911]==1) 
	 		intermediate[4095+2911:0+2911] <= intermediate[4095+2911:0+2911] + a; end
12'd2912: begin if(a[2912]==1) 
	 		intermediate[4095+2912:0+2912] <= intermediate[4095+2912:0+2912] + a; end
12'd2913: begin if(a[2913]==1) 
	 		intermediate[4095+2913:0+2913] <= intermediate[4095+2913:0+2913] + a; end
12'd2914: begin if(a[2914]==1) 
	 		intermediate[4095+2914:0+2914] <= intermediate[4095+2914:0+2914] + a; end
12'd2915: begin if(a[2915]==1) 
	 		intermediate[4095+2915:0+2915] <= intermediate[4095+2915:0+2915] + a; end
12'd2916: begin if(a[2916]==1) 
	 		intermediate[4095+2916:0+2916] <= intermediate[4095+2916:0+2916] + a; end
12'd2917: begin if(a[2917]==1) 
	 		intermediate[4095+2917:0+2917] <= intermediate[4095+2917:0+2917] + a; end
12'd2918: begin if(a[2918]==1) 
	 		intermediate[4095+2918:0+2918] <= intermediate[4095+2918:0+2918] + a; end
12'd2919: begin if(a[2919]==1) 
	 		intermediate[4095+2919:0+2919] <= intermediate[4095+2919:0+2919] + a; end
12'd2920: begin if(a[2920]==1) 
	 		intermediate[4095+2920:0+2920] <= intermediate[4095+2920:0+2920] + a; end
12'd2921: begin if(a[2921]==1) 
	 		intermediate[4095+2921:0+2921] <= intermediate[4095+2921:0+2921] + a; end
12'd2922: begin if(a[2922]==1) 
	 		intermediate[4095+2922:0+2922] <= intermediate[4095+2922:0+2922] + a; end
12'd2923: begin if(a[2923]==1) 
	 		intermediate[4095+2923:0+2923] <= intermediate[4095+2923:0+2923] + a; end
12'd2924: begin if(a[2924]==1) 
	 		intermediate[4095+2924:0+2924] <= intermediate[4095+2924:0+2924] + a; end
12'd2925: begin if(a[2925]==1) 
	 		intermediate[4095+2925:0+2925] <= intermediate[4095+2925:0+2925] + a; end
12'd2926: begin if(a[2926]==1) 
	 		intermediate[4095+2926:0+2926] <= intermediate[4095+2926:0+2926] + a; end
12'd2927: begin if(a[2927]==1) 
	 		intermediate[4095+2927:0+2927] <= intermediate[4095+2927:0+2927] + a; end
12'd2928: begin if(a[2928]==1) 
	 		intermediate[4095+2928:0+2928] <= intermediate[4095+2928:0+2928] + a; end
12'd2929: begin if(a[2929]==1) 
	 		intermediate[4095+2929:0+2929] <= intermediate[4095+2929:0+2929] + a; end
12'd2930: begin if(a[2930]==1) 
	 		intermediate[4095+2930:0+2930] <= intermediate[4095+2930:0+2930] + a; end
12'd2931: begin if(a[2931]==1) 
	 		intermediate[4095+2931:0+2931] <= intermediate[4095+2931:0+2931] + a; end
12'd2932: begin if(a[2932]==1) 
	 		intermediate[4095+2932:0+2932] <= intermediate[4095+2932:0+2932] + a; end
12'd2933: begin if(a[2933]==1) 
	 		intermediate[4095+2933:0+2933] <= intermediate[4095+2933:0+2933] + a; end
12'd2934: begin if(a[2934]==1) 
	 		intermediate[4095+2934:0+2934] <= intermediate[4095+2934:0+2934] + a; end
12'd2935: begin if(a[2935]==1) 
	 		intermediate[4095+2935:0+2935] <= intermediate[4095+2935:0+2935] + a; end
12'd2936: begin if(a[2936]==1) 
	 		intermediate[4095+2936:0+2936] <= intermediate[4095+2936:0+2936] + a; end
12'd2937: begin if(a[2937]==1) 
	 		intermediate[4095+2937:0+2937] <= intermediate[4095+2937:0+2937] + a; end
12'd2938: begin if(a[2938]==1) 
	 		intermediate[4095+2938:0+2938] <= intermediate[4095+2938:0+2938] + a; end
12'd2939: begin if(a[2939]==1) 
	 		intermediate[4095+2939:0+2939] <= intermediate[4095+2939:0+2939] + a; end
12'd2940: begin if(a[2940]==1) 
	 		intermediate[4095+2940:0+2940] <= intermediate[4095+2940:0+2940] + a; end
12'd2941: begin if(a[2941]==1) 
	 		intermediate[4095+2941:0+2941] <= intermediate[4095+2941:0+2941] + a; end
12'd2942: begin if(a[2942]==1) 
	 		intermediate[4095+2942:0+2942] <= intermediate[4095+2942:0+2942] + a; end
12'd2943: begin if(a[2943]==1) 
	 		intermediate[4095+2943:0+2943] <= intermediate[4095+2943:0+2943] + a; end
12'd2944: begin if(a[2944]==1) 
	 		intermediate[4095+2944:0+2944] <= intermediate[4095+2944:0+2944] + a; end
12'd2945: begin if(a[2945]==1) 
	 		intermediate[4095+2945:0+2945] <= intermediate[4095+2945:0+2945] + a; end
12'd2946: begin if(a[2946]==1) 
	 		intermediate[4095+2946:0+2946] <= intermediate[4095+2946:0+2946] + a; end
12'd2947: begin if(a[2947]==1) 
	 		intermediate[4095+2947:0+2947] <= intermediate[4095+2947:0+2947] + a; end
12'd2948: begin if(a[2948]==1) 
	 		intermediate[4095+2948:0+2948] <= intermediate[4095+2948:0+2948] + a; end
12'd2949: begin if(a[2949]==1) 
	 		intermediate[4095+2949:0+2949] <= intermediate[4095+2949:0+2949] + a; end
12'd2950: begin if(a[2950]==1) 
	 		intermediate[4095+2950:0+2950] <= intermediate[4095+2950:0+2950] + a; end
12'd2951: begin if(a[2951]==1) 
	 		intermediate[4095+2951:0+2951] <= intermediate[4095+2951:0+2951] + a; end
12'd2952: begin if(a[2952]==1) 
	 		intermediate[4095+2952:0+2952] <= intermediate[4095+2952:0+2952] + a; end
12'd2953: begin if(a[2953]==1) 
	 		intermediate[4095+2953:0+2953] <= intermediate[4095+2953:0+2953] + a; end
12'd2954: begin if(a[2954]==1) 
	 		intermediate[4095+2954:0+2954] <= intermediate[4095+2954:0+2954] + a; end
12'd2955: begin if(a[2955]==1) 
	 		intermediate[4095+2955:0+2955] <= intermediate[4095+2955:0+2955] + a; end
12'd2956: begin if(a[2956]==1) 
	 		intermediate[4095+2956:0+2956] <= intermediate[4095+2956:0+2956] + a; end
12'd2957: begin if(a[2957]==1) 
	 		intermediate[4095+2957:0+2957] <= intermediate[4095+2957:0+2957] + a; end
12'd2958: begin if(a[2958]==1) 
	 		intermediate[4095+2958:0+2958] <= intermediate[4095+2958:0+2958] + a; end
12'd2959: begin if(a[2959]==1) 
	 		intermediate[4095+2959:0+2959] <= intermediate[4095+2959:0+2959] + a; end
12'd2960: begin if(a[2960]==1) 
	 		intermediate[4095+2960:0+2960] <= intermediate[4095+2960:0+2960] + a; end
12'd2961: begin if(a[2961]==1) 
	 		intermediate[4095+2961:0+2961] <= intermediate[4095+2961:0+2961] + a; end
12'd2962: begin if(a[2962]==1) 
	 		intermediate[4095+2962:0+2962] <= intermediate[4095+2962:0+2962] + a; end
12'd2963: begin if(a[2963]==1) 
	 		intermediate[4095+2963:0+2963] <= intermediate[4095+2963:0+2963] + a; end
12'd2964: begin if(a[2964]==1) 
	 		intermediate[4095+2964:0+2964] <= intermediate[4095+2964:0+2964] + a; end
12'd2965: begin if(a[2965]==1) 
	 		intermediate[4095+2965:0+2965] <= intermediate[4095+2965:0+2965] + a; end
12'd2966: begin if(a[2966]==1) 
	 		intermediate[4095+2966:0+2966] <= intermediate[4095+2966:0+2966] + a; end
12'd2967: begin if(a[2967]==1) 
	 		intermediate[4095+2967:0+2967] <= intermediate[4095+2967:0+2967] + a; end
12'd2968: begin if(a[2968]==1) 
	 		intermediate[4095+2968:0+2968] <= intermediate[4095+2968:0+2968] + a; end
12'd2969: begin if(a[2969]==1) 
	 		intermediate[4095+2969:0+2969] <= intermediate[4095+2969:0+2969] + a; end
12'd2970: begin if(a[2970]==1) 
	 		intermediate[4095+2970:0+2970] <= intermediate[4095+2970:0+2970] + a; end
12'd2971: begin if(a[2971]==1) 
	 		intermediate[4095+2971:0+2971] <= intermediate[4095+2971:0+2971] + a; end
12'd2972: begin if(a[2972]==1) 
	 		intermediate[4095+2972:0+2972] <= intermediate[4095+2972:0+2972] + a; end
12'd2973: begin if(a[2973]==1) 
	 		intermediate[4095+2973:0+2973] <= intermediate[4095+2973:0+2973] + a; end
12'd2974: begin if(a[2974]==1) 
	 		intermediate[4095+2974:0+2974] <= intermediate[4095+2974:0+2974] + a; end
12'd2975: begin if(a[2975]==1) 
	 		intermediate[4095+2975:0+2975] <= intermediate[4095+2975:0+2975] + a; end
12'd2976: begin if(a[2976]==1) 
	 		intermediate[4095+2976:0+2976] <= intermediate[4095+2976:0+2976] + a; end
12'd2977: begin if(a[2977]==1) 
	 		intermediate[4095+2977:0+2977] <= intermediate[4095+2977:0+2977] + a; end
12'd2978: begin if(a[2978]==1) 
	 		intermediate[4095+2978:0+2978] <= intermediate[4095+2978:0+2978] + a; end
12'd2979: begin if(a[2979]==1) 
	 		intermediate[4095+2979:0+2979] <= intermediate[4095+2979:0+2979] + a; end
12'd2980: begin if(a[2980]==1) 
	 		intermediate[4095+2980:0+2980] <= intermediate[4095+2980:0+2980] + a; end
12'd2981: begin if(a[2981]==1) 
	 		intermediate[4095+2981:0+2981] <= intermediate[4095+2981:0+2981] + a; end
12'd2982: begin if(a[2982]==1) 
	 		intermediate[4095+2982:0+2982] <= intermediate[4095+2982:0+2982] + a; end
12'd2983: begin if(a[2983]==1) 
	 		intermediate[4095+2983:0+2983] <= intermediate[4095+2983:0+2983] + a; end
12'd2984: begin if(a[2984]==1) 
	 		intermediate[4095+2984:0+2984] <= intermediate[4095+2984:0+2984] + a; end
12'd2985: begin if(a[2985]==1) 
	 		intermediate[4095+2985:0+2985] <= intermediate[4095+2985:0+2985] + a; end
12'd2986: begin if(a[2986]==1) 
	 		intermediate[4095+2986:0+2986] <= intermediate[4095+2986:0+2986] + a; end
12'd2987: begin if(a[2987]==1) 
	 		intermediate[4095+2987:0+2987] <= intermediate[4095+2987:0+2987] + a; end
12'd2988: begin if(a[2988]==1) 
	 		intermediate[4095+2988:0+2988] <= intermediate[4095+2988:0+2988] + a; end
12'd2989: begin if(a[2989]==1) 
	 		intermediate[4095+2989:0+2989] <= intermediate[4095+2989:0+2989] + a; end
12'd2990: begin if(a[2990]==1) 
	 		intermediate[4095+2990:0+2990] <= intermediate[4095+2990:0+2990] + a; end
12'd2991: begin if(a[2991]==1) 
	 		intermediate[4095+2991:0+2991] <= intermediate[4095+2991:0+2991] + a; end
12'd2992: begin if(a[2992]==1) 
	 		intermediate[4095+2992:0+2992] <= intermediate[4095+2992:0+2992] + a; end
12'd2993: begin if(a[2993]==1) 
	 		intermediate[4095+2993:0+2993] <= intermediate[4095+2993:0+2993] + a; end
12'd2994: begin if(a[2994]==1) 
	 		intermediate[4095+2994:0+2994] <= intermediate[4095+2994:0+2994] + a; end
12'd2995: begin if(a[2995]==1) 
	 		intermediate[4095+2995:0+2995] <= intermediate[4095+2995:0+2995] + a; end
12'd2996: begin if(a[2996]==1) 
	 		intermediate[4095+2996:0+2996] <= intermediate[4095+2996:0+2996] + a; end
12'd2997: begin if(a[2997]==1) 
	 		intermediate[4095+2997:0+2997] <= intermediate[4095+2997:0+2997] + a; end
12'd2998: begin if(a[2998]==1) 
	 		intermediate[4095+2998:0+2998] <= intermediate[4095+2998:0+2998] + a; end
12'd2999: begin if(a[2999]==1) 
	 		intermediate[4095+2999:0+2999] <= intermediate[4095+2999:0+2999] + a; end
12'd3000: begin if(a[3000]==1) 
	 		intermediate[4095+3000:0+3000] <= intermediate[4095+3000:0+3000] + a; end
12'd3001: begin if(a[3001]==1) 
	 		intermediate[4095+3001:0+3001] <= intermediate[4095+3001:0+3001] + a; end
12'd3002: begin if(a[3002]==1) 
	 		intermediate[4095+3002:0+3002] <= intermediate[4095+3002:0+3002] + a; end
12'd3003: begin if(a[3003]==1) 
	 		intermediate[4095+3003:0+3003] <= intermediate[4095+3003:0+3003] + a; end
12'd3004: begin if(a[3004]==1) 
	 		intermediate[4095+3004:0+3004] <= intermediate[4095+3004:0+3004] + a; end
12'd3005: begin if(a[3005]==1) 
	 		intermediate[4095+3005:0+3005] <= intermediate[4095+3005:0+3005] + a; end
12'd3006: begin if(a[3006]==1) 
	 		intermediate[4095+3006:0+3006] <= intermediate[4095+3006:0+3006] + a; end
12'd3007: begin if(a[3007]==1) 
	 		intermediate[4095+3007:0+3007] <= intermediate[4095+3007:0+3007] + a; end
12'd3008: begin if(a[3008]==1) 
	 		intermediate[4095+3008:0+3008] <= intermediate[4095+3008:0+3008] + a; end
12'd3009: begin if(a[3009]==1) 
	 		intermediate[4095+3009:0+3009] <= intermediate[4095+3009:0+3009] + a; end
12'd3010: begin if(a[3010]==1) 
	 		intermediate[4095+3010:0+3010] <= intermediate[4095+3010:0+3010] + a; end
12'd3011: begin if(a[3011]==1) 
	 		intermediate[4095+3011:0+3011] <= intermediate[4095+3011:0+3011] + a; end
12'd3012: begin if(a[3012]==1) 
	 		intermediate[4095+3012:0+3012] <= intermediate[4095+3012:0+3012] + a; end
12'd3013: begin if(a[3013]==1) 
	 		intermediate[4095+3013:0+3013] <= intermediate[4095+3013:0+3013] + a; end
12'd3014: begin if(a[3014]==1) 
	 		intermediate[4095+3014:0+3014] <= intermediate[4095+3014:0+3014] + a; end
12'd3015: begin if(a[3015]==1) 
	 		intermediate[4095+3015:0+3015] <= intermediate[4095+3015:0+3015] + a; end
12'd3016: begin if(a[3016]==1) 
	 		intermediate[4095+3016:0+3016] <= intermediate[4095+3016:0+3016] + a; end
12'd3017: begin if(a[3017]==1) 
	 		intermediate[4095+3017:0+3017] <= intermediate[4095+3017:0+3017] + a; end
12'd3018: begin if(a[3018]==1) 
	 		intermediate[4095+3018:0+3018] <= intermediate[4095+3018:0+3018] + a; end
12'd3019: begin if(a[3019]==1) 
	 		intermediate[4095+3019:0+3019] <= intermediate[4095+3019:0+3019] + a; end
12'd3020: begin if(a[3020]==1) 
	 		intermediate[4095+3020:0+3020] <= intermediate[4095+3020:0+3020] + a; end
12'd3021: begin if(a[3021]==1) 
	 		intermediate[4095+3021:0+3021] <= intermediate[4095+3021:0+3021] + a; end
12'd3022: begin if(a[3022]==1) 
	 		intermediate[4095+3022:0+3022] <= intermediate[4095+3022:0+3022] + a; end
12'd3023: begin if(a[3023]==1) 
	 		intermediate[4095+3023:0+3023] <= intermediate[4095+3023:0+3023] + a; end
12'd3024: begin if(a[3024]==1) 
	 		intermediate[4095+3024:0+3024] <= intermediate[4095+3024:0+3024] + a; end
12'd3025: begin if(a[3025]==1) 
	 		intermediate[4095+3025:0+3025] <= intermediate[4095+3025:0+3025] + a; end
12'd3026: begin if(a[3026]==1) 
	 		intermediate[4095+3026:0+3026] <= intermediate[4095+3026:0+3026] + a; end
12'd3027: begin if(a[3027]==1) 
	 		intermediate[4095+3027:0+3027] <= intermediate[4095+3027:0+3027] + a; end
12'd3028: begin if(a[3028]==1) 
	 		intermediate[4095+3028:0+3028] <= intermediate[4095+3028:0+3028] + a; end
12'd3029: begin if(a[3029]==1) 
	 		intermediate[4095+3029:0+3029] <= intermediate[4095+3029:0+3029] + a; end
12'd3030: begin if(a[3030]==1) 
	 		intermediate[4095+3030:0+3030] <= intermediate[4095+3030:0+3030] + a; end
12'd3031: begin if(a[3031]==1) 
	 		intermediate[4095+3031:0+3031] <= intermediate[4095+3031:0+3031] + a; end
12'd3032: begin if(a[3032]==1) 
	 		intermediate[4095+3032:0+3032] <= intermediate[4095+3032:0+3032] + a; end
12'd3033: begin if(a[3033]==1) 
	 		intermediate[4095+3033:0+3033] <= intermediate[4095+3033:0+3033] + a; end
12'd3034: begin if(a[3034]==1) 
	 		intermediate[4095+3034:0+3034] <= intermediate[4095+3034:0+3034] + a; end
12'd3035: begin if(a[3035]==1) 
	 		intermediate[4095+3035:0+3035] <= intermediate[4095+3035:0+3035] + a; end
12'd3036: begin if(a[3036]==1) 
	 		intermediate[4095+3036:0+3036] <= intermediate[4095+3036:0+3036] + a; end
12'd3037: begin if(a[3037]==1) 
	 		intermediate[4095+3037:0+3037] <= intermediate[4095+3037:0+3037] + a; end
12'd3038: begin if(a[3038]==1) 
	 		intermediate[4095+3038:0+3038] <= intermediate[4095+3038:0+3038] + a; end
12'd3039: begin if(a[3039]==1) 
	 		intermediate[4095+3039:0+3039] <= intermediate[4095+3039:0+3039] + a; end
12'd3040: begin if(a[3040]==1) 
	 		intermediate[4095+3040:0+3040] <= intermediate[4095+3040:0+3040] + a; end
12'd3041: begin if(a[3041]==1) 
	 		intermediate[4095+3041:0+3041] <= intermediate[4095+3041:0+3041] + a; end
12'd3042: begin if(a[3042]==1) 
	 		intermediate[4095+3042:0+3042] <= intermediate[4095+3042:0+3042] + a; end
12'd3043: begin if(a[3043]==1) 
	 		intermediate[4095+3043:0+3043] <= intermediate[4095+3043:0+3043] + a; end
12'd3044: begin if(a[3044]==1) 
	 		intermediate[4095+3044:0+3044] <= intermediate[4095+3044:0+3044] + a; end
12'd3045: begin if(a[3045]==1) 
	 		intermediate[4095+3045:0+3045] <= intermediate[4095+3045:0+3045] + a; end
12'd3046: begin if(a[3046]==1) 
	 		intermediate[4095+3046:0+3046] <= intermediate[4095+3046:0+3046] + a; end
12'd3047: begin if(a[3047]==1) 
	 		intermediate[4095+3047:0+3047] <= intermediate[4095+3047:0+3047] + a; end
12'd3048: begin if(a[3048]==1) 
	 		intermediate[4095+3048:0+3048] <= intermediate[4095+3048:0+3048] + a; end
12'd3049: begin if(a[3049]==1) 
	 		intermediate[4095+3049:0+3049] <= intermediate[4095+3049:0+3049] + a; end
12'd3050: begin if(a[3050]==1) 
	 		intermediate[4095+3050:0+3050] <= intermediate[4095+3050:0+3050] + a; end
12'd3051: begin if(a[3051]==1) 
	 		intermediate[4095+3051:0+3051] <= intermediate[4095+3051:0+3051] + a; end
12'd3052: begin if(a[3052]==1) 
	 		intermediate[4095+3052:0+3052] <= intermediate[4095+3052:0+3052] + a; end
12'd3053: begin if(a[3053]==1) 
	 		intermediate[4095+3053:0+3053] <= intermediate[4095+3053:0+3053] + a; end
12'd3054: begin if(a[3054]==1) 
	 		intermediate[4095+3054:0+3054] <= intermediate[4095+3054:0+3054] + a; end
12'd3055: begin if(a[3055]==1) 
	 		intermediate[4095+3055:0+3055] <= intermediate[4095+3055:0+3055] + a; end
12'd3056: begin if(a[3056]==1) 
	 		intermediate[4095+3056:0+3056] <= intermediate[4095+3056:0+3056] + a; end
12'd3057: begin if(a[3057]==1) 
	 		intermediate[4095+3057:0+3057] <= intermediate[4095+3057:0+3057] + a; end
12'd3058: begin if(a[3058]==1) 
	 		intermediate[4095+3058:0+3058] <= intermediate[4095+3058:0+3058] + a; end
12'd3059: begin if(a[3059]==1) 
	 		intermediate[4095+3059:0+3059] <= intermediate[4095+3059:0+3059] + a; end
12'd3060: begin if(a[3060]==1) 
	 		intermediate[4095+3060:0+3060] <= intermediate[4095+3060:0+3060] + a; end
12'd3061: begin if(a[3061]==1) 
	 		intermediate[4095+3061:0+3061] <= intermediate[4095+3061:0+3061] + a; end
12'd3062: begin if(a[3062]==1) 
	 		intermediate[4095+3062:0+3062] <= intermediate[4095+3062:0+3062] + a; end
12'd3063: begin if(a[3063]==1) 
	 		intermediate[4095+3063:0+3063] <= intermediate[4095+3063:0+3063] + a; end
12'd3064: begin if(a[3064]==1) 
	 		intermediate[4095+3064:0+3064] <= intermediate[4095+3064:0+3064] + a; end
12'd3065: begin if(a[3065]==1) 
	 		intermediate[4095+3065:0+3065] <= intermediate[4095+3065:0+3065] + a; end
12'd3066: begin if(a[3066]==1) 
	 		intermediate[4095+3066:0+3066] <= intermediate[4095+3066:0+3066] + a; end
12'd3067: begin if(a[3067]==1) 
	 		intermediate[4095+3067:0+3067] <= intermediate[4095+3067:0+3067] + a; end
12'd3068: begin if(a[3068]==1) 
	 		intermediate[4095+3068:0+3068] <= intermediate[4095+3068:0+3068] + a; end
12'd3069: begin if(a[3069]==1) 
	 		intermediate[4095+3069:0+3069] <= intermediate[4095+3069:0+3069] + a; end
12'd3070: begin if(a[3070]==1) 
	 		intermediate[4095+3070:0+3070] <= intermediate[4095+3070:0+3070] + a; end
12'd3071: begin if(a[3071]==1) 
	 		intermediate[4095+3071:0+3071] <= intermediate[4095+3071:0+3071] + a; end
12'd3072: begin if(a[3072]==1) 
	 		intermediate[4095+3072:0+3072] <= intermediate[4095+3072:0+3072] + a; end
12'd3073: begin if(a[3073]==1) 
	 		intermediate[4095+3073:0+3073] <= intermediate[4095+3073:0+3073] + a; end
12'd3074: begin if(a[3074]==1) 
	 		intermediate[4095+3074:0+3074] <= intermediate[4095+3074:0+3074] + a; end
12'd3075: begin if(a[3075]==1) 
	 		intermediate[4095+3075:0+3075] <= intermediate[4095+3075:0+3075] + a; end
12'd3076: begin if(a[3076]==1) 
	 		intermediate[4095+3076:0+3076] <= intermediate[4095+3076:0+3076] + a; end
12'd3077: begin if(a[3077]==1) 
	 		intermediate[4095+3077:0+3077] <= intermediate[4095+3077:0+3077] + a; end
12'd3078: begin if(a[3078]==1) 
	 		intermediate[4095+3078:0+3078] <= intermediate[4095+3078:0+3078] + a; end
12'd3079: begin if(a[3079]==1) 
	 		intermediate[4095+3079:0+3079] <= intermediate[4095+3079:0+3079] + a; end
12'd3080: begin if(a[3080]==1) 
	 		intermediate[4095+3080:0+3080] <= intermediate[4095+3080:0+3080] + a; end
12'd3081: begin if(a[3081]==1) 
	 		intermediate[4095+3081:0+3081] <= intermediate[4095+3081:0+3081] + a; end
12'd3082: begin if(a[3082]==1) 
	 		intermediate[4095+3082:0+3082] <= intermediate[4095+3082:0+3082] + a; end
12'd3083: begin if(a[3083]==1) 
	 		intermediate[4095+3083:0+3083] <= intermediate[4095+3083:0+3083] + a; end
12'd3084: begin if(a[3084]==1) 
	 		intermediate[4095+3084:0+3084] <= intermediate[4095+3084:0+3084] + a; end
12'd3085: begin if(a[3085]==1) 
	 		intermediate[4095+3085:0+3085] <= intermediate[4095+3085:0+3085] + a; end
12'd3086: begin if(a[3086]==1) 
	 		intermediate[4095+3086:0+3086] <= intermediate[4095+3086:0+3086] + a; end
12'd3087: begin if(a[3087]==1) 
	 		intermediate[4095+3087:0+3087] <= intermediate[4095+3087:0+3087] + a; end
12'd3088: begin if(a[3088]==1) 
	 		intermediate[4095+3088:0+3088] <= intermediate[4095+3088:0+3088] + a; end
12'd3089: begin if(a[3089]==1) 
	 		intermediate[4095+3089:0+3089] <= intermediate[4095+3089:0+3089] + a; end
12'd3090: begin if(a[3090]==1) 
	 		intermediate[4095+3090:0+3090] <= intermediate[4095+3090:0+3090] + a; end
12'd3091: begin if(a[3091]==1) 
	 		intermediate[4095+3091:0+3091] <= intermediate[4095+3091:0+3091] + a; end
12'd3092: begin if(a[3092]==1) 
	 		intermediate[4095+3092:0+3092] <= intermediate[4095+3092:0+3092] + a; end
12'd3093: begin if(a[3093]==1) 
	 		intermediate[4095+3093:0+3093] <= intermediate[4095+3093:0+3093] + a; end
12'd3094: begin if(a[3094]==1) 
	 		intermediate[4095+3094:0+3094] <= intermediate[4095+3094:0+3094] + a; end
12'd3095: begin if(a[3095]==1) 
	 		intermediate[4095+3095:0+3095] <= intermediate[4095+3095:0+3095] + a; end
12'd3096: begin if(a[3096]==1) 
	 		intermediate[4095+3096:0+3096] <= intermediate[4095+3096:0+3096] + a; end
12'd3097: begin if(a[3097]==1) 
	 		intermediate[4095+3097:0+3097] <= intermediate[4095+3097:0+3097] + a; end
12'd3098: begin if(a[3098]==1) 
	 		intermediate[4095+3098:0+3098] <= intermediate[4095+3098:0+3098] + a; end
12'd3099: begin if(a[3099]==1) 
	 		intermediate[4095+3099:0+3099] <= intermediate[4095+3099:0+3099] + a; end
12'd3100: begin if(a[3100]==1) 
	 		intermediate[4095+3100:0+3100] <= intermediate[4095+3100:0+3100] + a; end
12'd3101: begin if(a[3101]==1) 
	 		intermediate[4095+3101:0+3101] <= intermediate[4095+3101:0+3101] + a; end
12'd3102: begin if(a[3102]==1) 
	 		intermediate[4095+3102:0+3102] <= intermediate[4095+3102:0+3102] + a; end
12'd3103: begin if(a[3103]==1) 
	 		intermediate[4095+3103:0+3103] <= intermediate[4095+3103:0+3103] + a; end
12'd3104: begin if(a[3104]==1) 
	 		intermediate[4095+3104:0+3104] <= intermediate[4095+3104:0+3104] + a; end
12'd3105: begin if(a[3105]==1) 
	 		intermediate[4095+3105:0+3105] <= intermediate[4095+3105:0+3105] + a; end
12'd3106: begin if(a[3106]==1) 
	 		intermediate[4095+3106:0+3106] <= intermediate[4095+3106:0+3106] + a; end
12'd3107: begin if(a[3107]==1) 
	 		intermediate[4095+3107:0+3107] <= intermediate[4095+3107:0+3107] + a; end
12'd3108: begin if(a[3108]==1) 
	 		intermediate[4095+3108:0+3108] <= intermediate[4095+3108:0+3108] + a; end
12'd3109: begin if(a[3109]==1) 
	 		intermediate[4095+3109:0+3109] <= intermediate[4095+3109:0+3109] + a; end
12'd3110: begin if(a[3110]==1) 
	 		intermediate[4095+3110:0+3110] <= intermediate[4095+3110:0+3110] + a; end
12'd3111: begin if(a[3111]==1) 
	 		intermediate[4095+3111:0+3111] <= intermediate[4095+3111:0+3111] + a; end
12'd3112: begin if(a[3112]==1) 
	 		intermediate[4095+3112:0+3112] <= intermediate[4095+3112:0+3112] + a; end
12'd3113: begin if(a[3113]==1) 
	 		intermediate[4095+3113:0+3113] <= intermediate[4095+3113:0+3113] + a; end
12'd3114: begin if(a[3114]==1) 
	 		intermediate[4095+3114:0+3114] <= intermediate[4095+3114:0+3114] + a; end
12'd3115: begin if(a[3115]==1) 
	 		intermediate[4095+3115:0+3115] <= intermediate[4095+3115:0+3115] + a; end
12'd3116: begin if(a[3116]==1) 
	 		intermediate[4095+3116:0+3116] <= intermediate[4095+3116:0+3116] + a; end
12'd3117: begin if(a[3117]==1) 
	 		intermediate[4095+3117:0+3117] <= intermediate[4095+3117:0+3117] + a; end
12'd3118: begin if(a[3118]==1) 
	 		intermediate[4095+3118:0+3118] <= intermediate[4095+3118:0+3118] + a; end
12'd3119: begin if(a[3119]==1) 
	 		intermediate[4095+3119:0+3119] <= intermediate[4095+3119:0+3119] + a; end
12'd3120: begin if(a[3120]==1) 
	 		intermediate[4095+3120:0+3120] <= intermediate[4095+3120:0+3120] + a; end
12'd3121: begin if(a[3121]==1) 
	 		intermediate[4095+3121:0+3121] <= intermediate[4095+3121:0+3121] + a; end
12'd3122: begin if(a[3122]==1) 
	 		intermediate[4095+3122:0+3122] <= intermediate[4095+3122:0+3122] + a; end
12'd3123: begin if(a[3123]==1) 
	 		intermediate[4095+3123:0+3123] <= intermediate[4095+3123:0+3123] + a; end
12'd3124: begin if(a[3124]==1) 
	 		intermediate[4095+3124:0+3124] <= intermediate[4095+3124:0+3124] + a; end
12'd3125: begin if(a[3125]==1) 
	 		intermediate[4095+3125:0+3125] <= intermediate[4095+3125:0+3125] + a; end
12'd3126: begin if(a[3126]==1) 
	 		intermediate[4095+3126:0+3126] <= intermediate[4095+3126:0+3126] + a; end
12'd3127: begin if(a[3127]==1) 
	 		intermediate[4095+3127:0+3127] <= intermediate[4095+3127:0+3127] + a; end
12'd3128: begin if(a[3128]==1) 
	 		intermediate[4095+3128:0+3128] <= intermediate[4095+3128:0+3128] + a; end
12'd3129: begin if(a[3129]==1) 
	 		intermediate[4095+3129:0+3129] <= intermediate[4095+3129:0+3129] + a; end
12'd3130: begin if(a[3130]==1) 
	 		intermediate[4095+3130:0+3130] <= intermediate[4095+3130:0+3130] + a; end
12'd3131: begin if(a[3131]==1) 
	 		intermediate[4095+3131:0+3131] <= intermediate[4095+3131:0+3131] + a; end
12'd3132: begin if(a[3132]==1) 
	 		intermediate[4095+3132:0+3132] <= intermediate[4095+3132:0+3132] + a; end
12'd3133: begin if(a[3133]==1) 
	 		intermediate[4095+3133:0+3133] <= intermediate[4095+3133:0+3133] + a; end
12'd3134: begin if(a[3134]==1) 
	 		intermediate[4095+3134:0+3134] <= intermediate[4095+3134:0+3134] + a; end
12'd3135: begin if(a[3135]==1) 
	 		intermediate[4095+3135:0+3135] <= intermediate[4095+3135:0+3135] + a; end
12'd3136: begin if(a[3136]==1) 
	 		intermediate[4095+3136:0+3136] <= intermediate[4095+3136:0+3136] + a; end
12'd3137: begin if(a[3137]==1) 
	 		intermediate[4095+3137:0+3137] <= intermediate[4095+3137:0+3137] + a; end
12'd3138: begin if(a[3138]==1) 
	 		intermediate[4095+3138:0+3138] <= intermediate[4095+3138:0+3138] + a; end
12'd3139: begin if(a[3139]==1) 
	 		intermediate[4095+3139:0+3139] <= intermediate[4095+3139:0+3139] + a; end
12'd3140: begin if(a[3140]==1) 
	 		intermediate[4095+3140:0+3140] <= intermediate[4095+3140:0+3140] + a; end
12'd3141: begin if(a[3141]==1) 
	 		intermediate[4095+3141:0+3141] <= intermediate[4095+3141:0+3141] + a; end
12'd3142: begin if(a[3142]==1) 
	 		intermediate[4095+3142:0+3142] <= intermediate[4095+3142:0+3142] + a; end
12'd3143: begin if(a[3143]==1) 
	 		intermediate[4095+3143:0+3143] <= intermediate[4095+3143:0+3143] + a; end
12'd3144: begin if(a[3144]==1) 
	 		intermediate[4095+3144:0+3144] <= intermediate[4095+3144:0+3144] + a; end
12'd3145: begin if(a[3145]==1) 
	 		intermediate[4095+3145:0+3145] <= intermediate[4095+3145:0+3145] + a; end
12'd3146: begin if(a[3146]==1) 
	 		intermediate[4095+3146:0+3146] <= intermediate[4095+3146:0+3146] + a; end
12'd3147: begin if(a[3147]==1) 
	 		intermediate[4095+3147:0+3147] <= intermediate[4095+3147:0+3147] + a; end
12'd3148: begin if(a[3148]==1) 
	 		intermediate[4095+3148:0+3148] <= intermediate[4095+3148:0+3148] + a; end
12'd3149: begin if(a[3149]==1) 
	 		intermediate[4095+3149:0+3149] <= intermediate[4095+3149:0+3149] + a; end
12'd3150: begin if(a[3150]==1) 
	 		intermediate[4095+3150:0+3150] <= intermediate[4095+3150:0+3150] + a; end
12'd3151: begin if(a[3151]==1) 
	 		intermediate[4095+3151:0+3151] <= intermediate[4095+3151:0+3151] + a; end
12'd3152: begin if(a[3152]==1) 
	 		intermediate[4095+3152:0+3152] <= intermediate[4095+3152:0+3152] + a; end
12'd3153: begin if(a[3153]==1) 
	 		intermediate[4095+3153:0+3153] <= intermediate[4095+3153:0+3153] + a; end
12'd3154: begin if(a[3154]==1) 
	 		intermediate[4095+3154:0+3154] <= intermediate[4095+3154:0+3154] + a; end
12'd3155: begin if(a[3155]==1) 
	 		intermediate[4095+3155:0+3155] <= intermediate[4095+3155:0+3155] + a; end
12'd3156: begin if(a[3156]==1) 
	 		intermediate[4095+3156:0+3156] <= intermediate[4095+3156:0+3156] + a; end
12'd3157: begin if(a[3157]==1) 
	 		intermediate[4095+3157:0+3157] <= intermediate[4095+3157:0+3157] + a; end
12'd3158: begin if(a[3158]==1) 
	 		intermediate[4095+3158:0+3158] <= intermediate[4095+3158:0+3158] + a; end
12'd3159: begin if(a[3159]==1) 
	 		intermediate[4095+3159:0+3159] <= intermediate[4095+3159:0+3159] + a; end
12'd3160: begin if(a[3160]==1) 
	 		intermediate[4095+3160:0+3160] <= intermediate[4095+3160:0+3160] + a; end
12'd3161: begin if(a[3161]==1) 
	 		intermediate[4095+3161:0+3161] <= intermediate[4095+3161:0+3161] + a; end
12'd3162: begin if(a[3162]==1) 
	 		intermediate[4095+3162:0+3162] <= intermediate[4095+3162:0+3162] + a; end
12'd3163: begin if(a[3163]==1) 
	 		intermediate[4095+3163:0+3163] <= intermediate[4095+3163:0+3163] + a; end
12'd3164: begin if(a[3164]==1) 
	 		intermediate[4095+3164:0+3164] <= intermediate[4095+3164:0+3164] + a; end
12'd3165: begin if(a[3165]==1) 
	 		intermediate[4095+3165:0+3165] <= intermediate[4095+3165:0+3165] + a; end
12'd3166: begin if(a[3166]==1) 
	 		intermediate[4095+3166:0+3166] <= intermediate[4095+3166:0+3166] + a; end
12'd3167: begin if(a[3167]==1) 
	 		intermediate[4095+3167:0+3167] <= intermediate[4095+3167:0+3167] + a; end
12'd3168: begin if(a[3168]==1) 
	 		intermediate[4095+3168:0+3168] <= intermediate[4095+3168:0+3168] + a; end
12'd3169: begin if(a[3169]==1) 
	 		intermediate[4095+3169:0+3169] <= intermediate[4095+3169:0+3169] + a; end
12'd3170: begin if(a[3170]==1) 
	 		intermediate[4095+3170:0+3170] <= intermediate[4095+3170:0+3170] + a; end
12'd3171: begin if(a[3171]==1) 
	 		intermediate[4095+3171:0+3171] <= intermediate[4095+3171:0+3171] + a; end
12'd3172: begin if(a[3172]==1) 
	 		intermediate[4095+3172:0+3172] <= intermediate[4095+3172:0+3172] + a; end
12'd3173: begin if(a[3173]==1) 
	 		intermediate[4095+3173:0+3173] <= intermediate[4095+3173:0+3173] + a; end
12'd3174: begin if(a[3174]==1) 
	 		intermediate[4095+3174:0+3174] <= intermediate[4095+3174:0+3174] + a; end
12'd3175: begin if(a[3175]==1) 
	 		intermediate[4095+3175:0+3175] <= intermediate[4095+3175:0+3175] + a; end
12'd3176: begin if(a[3176]==1) 
	 		intermediate[4095+3176:0+3176] <= intermediate[4095+3176:0+3176] + a; end
12'd3177: begin if(a[3177]==1) 
	 		intermediate[4095+3177:0+3177] <= intermediate[4095+3177:0+3177] + a; end
12'd3178: begin if(a[3178]==1) 
	 		intermediate[4095+3178:0+3178] <= intermediate[4095+3178:0+3178] + a; end
12'd3179: begin if(a[3179]==1) 
	 		intermediate[4095+3179:0+3179] <= intermediate[4095+3179:0+3179] + a; end
12'd3180: begin if(a[3180]==1) 
	 		intermediate[4095+3180:0+3180] <= intermediate[4095+3180:0+3180] + a; end
12'd3181: begin if(a[3181]==1) 
	 		intermediate[4095+3181:0+3181] <= intermediate[4095+3181:0+3181] + a; end
12'd3182: begin if(a[3182]==1) 
	 		intermediate[4095+3182:0+3182] <= intermediate[4095+3182:0+3182] + a; end
12'd3183: begin if(a[3183]==1) 
	 		intermediate[4095+3183:0+3183] <= intermediate[4095+3183:0+3183] + a; end
12'd3184: begin if(a[3184]==1) 
	 		intermediate[4095+3184:0+3184] <= intermediate[4095+3184:0+3184] + a; end
12'd3185: begin if(a[3185]==1) 
	 		intermediate[4095+3185:0+3185] <= intermediate[4095+3185:0+3185] + a; end
12'd3186: begin if(a[3186]==1) 
	 		intermediate[4095+3186:0+3186] <= intermediate[4095+3186:0+3186] + a; end
12'd3187: begin if(a[3187]==1) 
	 		intermediate[4095+3187:0+3187] <= intermediate[4095+3187:0+3187] + a; end
12'd3188: begin if(a[3188]==1) 
	 		intermediate[4095+3188:0+3188] <= intermediate[4095+3188:0+3188] + a; end
12'd3189: begin if(a[3189]==1) 
	 		intermediate[4095+3189:0+3189] <= intermediate[4095+3189:0+3189] + a; end
12'd3190: begin if(a[3190]==1) 
	 		intermediate[4095+3190:0+3190] <= intermediate[4095+3190:0+3190] + a; end
12'd3191: begin if(a[3191]==1) 
	 		intermediate[4095+3191:0+3191] <= intermediate[4095+3191:0+3191] + a; end
12'd3192: begin if(a[3192]==1) 
	 		intermediate[4095+3192:0+3192] <= intermediate[4095+3192:0+3192] + a; end
12'd3193: begin if(a[3193]==1) 
	 		intermediate[4095+3193:0+3193] <= intermediate[4095+3193:0+3193] + a; end
12'd3194: begin if(a[3194]==1) 
	 		intermediate[4095+3194:0+3194] <= intermediate[4095+3194:0+3194] + a; end
12'd3195: begin if(a[3195]==1) 
	 		intermediate[4095+3195:0+3195] <= intermediate[4095+3195:0+3195] + a; end
12'd3196: begin if(a[3196]==1) 
	 		intermediate[4095+3196:0+3196] <= intermediate[4095+3196:0+3196] + a; end
12'd3197: begin if(a[3197]==1) 
	 		intermediate[4095+3197:0+3197] <= intermediate[4095+3197:0+3197] + a; end
12'd3198: begin if(a[3198]==1) 
	 		intermediate[4095+3198:0+3198] <= intermediate[4095+3198:0+3198] + a; end
12'd3199: begin if(a[3199]==1) 
	 		intermediate[4095+3199:0+3199] <= intermediate[4095+3199:0+3199] + a; end
12'd3200: begin if(a[3200]==1) 
	 		intermediate[4095+3200:0+3200] <= intermediate[4095+3200:0+3200] + a; end
12'd3201: begin if(a[3201]==1) 
	 		intermediate[4095+3201:0+3201] <= intermediate[4095+3201:0+3201] + a; end
12'd3202: begin if(a[3202]==1) 
	 		intermediate[4095+3202:0+3202] <= intermediate[4095+3202:0+3202] + a; end
12'd3203: begin if(a[3203]==1) 
	 		intermediate[4095+3203:0+3203] <= intermediate[4095+3203:0+3203] + a; end
12'd3204: begin if(a[3204]==1) 
	 		intermediate[4095+3204:0+3204] <= intermediate[4095+3204:0+3204] + a; end
12'd3205: begin if(a[3205]==1) 
	 		intermediate[4095+3205:0+3205] <= intermediate[4095+3205:0+3205] + a; end
12'd3206: begin if(a[3206]==1) 
	 		intermediate[4095+3206:0+3206] <= intermediate[4095+3206:0+3206] + a; end
12'd3207: begin if(a[3207]==1) 
	 		intermediate[4095+3207:0+3207] <= intermediate[4095+3207:0+3207] + a; end
12'd3208: begin if(a[3208]==1) 
	 		intermediate[4095+3208:0+3208] <= intermediate[4095+3208:0+3208] + a; end
12'd3209: begin if(a[3209]==1) 
	 		intermediate[4095+3209:0+3209] <= intermediate[4095+3209:0+3209] + a; end
12'd3210: begin if(a[3210]==1) 
	 		intermediate[4095+3210:0+3210] <= intermediate[4095+3210:0+3210] + a; end
12'd3211: begin if(a[3211]==1) 
	 		intermediate[4095+3211:0+3211] <= intermediate[4095+3211:0+3211] + a; end
12'd3212: begin if(a[3212]==1) 
	 		intermediate[4095+3212:0+3212] <= intermediate[4095+3212:0+3212] + a; end
12'd3213: begin if(a[3213]==1) 
	 		intermediate[4095+3213:0+3213] <= intermediate[4095+3213:0+3213] + a; end
12'd3214: begin if(a[3214]==1) 
	 		intermediate[4095+3214:0+3214] <= intermediate[4095+3214:0+3214] + a; end
12'd3215: begin if(a[3215]==1) 
	 		intermediate[4095+3215:0+3215] <= intermediate[4095+3215:0+3215] + a; end
12'd3216: begin if(a[3216]==1) 
	 		intermediate[4095+3216:0+3216] <= intermediate[4095+3216:0+3216] + a; end
12'd3217: begin if(a[3217]==1) 
	 		intermediate[4095+3217:0+3217] <= intermediate[4095+3217:0+3217] + a; end
12'd3218: begin if(a[3218]==1) 
	 		intermediate[4095+3218:0+3218] <= intermediate[4095+3218:0+3218] + a; end
12'd3219: begin if(a[3219]==1) 
	 		intermediate[4095+3219:0+3219] <= intermediate[4095+3219:0+3219] + a; end
12'd3220: begin if(a[3220]==1) 
	 		intermediate[4095+3220:0+3220] <= intermediate[4095+3220:0+3220] + a; end
12'd3221: begin if(a[3221]==1) 
	 		intermediate[4095+3221:0+3221] <= intermediate[4095+3221:0+3221] + a; end
12'd3222: begin if(a[3222]==1) 
	 		intermediate[4095+3222:0+3222] <= intermediate[4095+3222:0+3222] + a; end
12'd3223: begin if(a[3223]==1) 
	 		intermediate[4095+3223:0+3223] <= intermediate[4095+3223:0+3223] + a; end
12'd3224: begin if(a[3224]==1) 
	 		intermediate[4095+3224:0+3224] <= intermediate[4095+3224:0+3224] + a; end
12'd3225: begin if(a[3225]==1) 
	 		intermediate[4095+3225:0+3225] <= intermediate[4095+3225:0+3225] + a; end
12'd3226: begin if(a[3226]==1) 
	 		intermediate[4095+3226:0+3226] <= intermediate[4095+3226:0+3226] + a; end
12'd3227: begin if(a[3227]==1) 
	 		intermediate[4095+3227:0+3227] <= intermediate[4095+3227:0+3227] + a; end
12'd3228: begin if(a[3228]==1) 
	 		intermediate[4095+3228:0+3228] <= intermediate[4095+3228:0+3228] + a; end
12'd3229: begin if(a[3229]==1) 
	 		intermediate[4095+3229:0+3229] <= intermediate[4095+3229:0+3229] + a; end
12'd3230: begin if(a[3230]==1) 
	 		intermediate[4095+3230:0+3230] <= intermediate[4095+3230:0+3230] + a; end
12'd3231: begin if(a[3231]==1) 
	 		intermediate[4095+3231:0+3231] <= intermediate[4095+3231:0+3231] + a; end
12'd3232: begin if(a[3232]==1) 
	 		intermediate[4095+3232:0+3232] <= intermediate[4095+3232:0+3232] + a; end
12'd3233: begin if(a[3233]==1) 
	 		intermediate[4095+3233:0+3233] <= intermediate[4095+3233:0+3233] + a; end
12'd3234: begin if(a[3234]==1) 
	 		intermediate[4095+3234:0+3234] <= intermediate[4095+3234:0+3234] + a; end
12'd3235: begin if(a[3235]==1) 
	 		intermediate[4095+3235:0+3235] <= intermediate[4095+3235:0+3235] + a; end
12'd3236: begin if(a[3236]==1) 
	 		intermediate[4095+3236:0+3236] <= intermediate[4095+3236:0+3236] + a; end
12'd3237: begin if(a[3237]==1) 
	 		intermediate[4095+3237:0+3237] <= intermediate[4095+3237:0+3237] + a; end
12'd3238: begin if(a[3238]==1) 
	 		intermediate[4095+3238:0+3238] <= intermediate[4095+3238:0+3238] + a; end
12'd3239: begin if(a[3239]==1) 
	 		intermediate[4095+3239:0+3239] <= intermediate[4095+3239:0+3239] + a; end
12'd3240: begin if(a[3240]==1) 
	 		intermediate[4095+3240:0+3240] <= intermediate[4095+3240:0+3240] + a; end
12'd3241: begin if(a[3241]==1) 
	 		intermediate[4095+3241:0+3241] <= intermediate[4095+3241:0+3241] + a; end
12'd3242: begin if(a[3242]==1) 
	 		intermediate[4095+3242:0+3242] <= intermediate[4095+3242:0+3242] + a; end
12'd3243: begin if(a[3243]==1) 
	 		intermediate[4095+3243:0+3243] <= intermediate[4095+3243:0+3243] + a; end
12'd3244: begin if(a[3244]==1) 
	 		intermediate[4095+3244:0+3244] <= intermediate[4095+3244:0+3244] + a; end
12'd3245: begin if(a[3245]==1) 
	 		intermediate[4095+3245:0+3245] <= intermediate[4095+3245:0+3245] + a; end
12'd3246: begin if(a[3246]==1) 
	 		intermediate[4095+3246:0+3246] <= intermediate[4095+3246:0+3246] + a; end
12'd3247: begin if(a[3247]==1) 
	 		intermediate[4095+3247:0+3247] <= intermediate[4095+3247:0+3247] + a; end
12'd3248: begin if(a[3248]==1) 
	 		intermediate[4095+3248:0+3248] <= intermediate[4095+3248:0+3248] + a; end
12'd3249: begin if(a[3249]==1) 
	 		intermediate[4095+3249:0+3249] <= intermediate[4095+3249:0+3249] + a; end
12'd3250: begin if(a[3250]==1) 
	 		intermediate[4095+3250:0+3250] <= intermediate[4095+3250:0+3250] + a; end
12'd3251: begin if(a[3251]==1) 
	 		intermediate[4095+3251:0+3251] <= intermediate[4095+3251:0+3251] + a; end
12'd3252: begin if(a[3252]==1) 
	 		intermediate[4095+3252:0+3252] <= intermediate[4095+3252:0+3252] + a; end
12'd3253: begin if(a[3253]==1) 
	 		intermediate[4095+3253:0+3253] <= intermediate[4095+3253:0+3253] + a; end
12'd3254: begin if(a[3254]==1) 
	 		intermediate[4095+3254:0+3254] <= intermediate[4095+3254:0+3254] + a; end
12'd3255: begin if(a[3255]==1) 
	 		intermediate[4095+3255:0+3255] <= intermediate[4095+3255:0+3255] + a; end
12'd3256: begin if(a[3256]==1) 
	 		intermediate[4095+3256:0+3256] <= intermediate[4095+3256:0+3256] + a; end
12'd3257: begin if(a[3257]==1) 
	 		intermediate[4095+3257:0+3257] <= intermediate[4095+3257:0+3257] + a; end
12'd3258: begin if(a[3258]==1) 
	 		intermediate[4095+3258:0+3258] <= intermediate[4095+3258:0+3258] + a; end
12'd3259: begin if(a[3259]==1) 
	 		intermediate[4095+3259:0+3259] <= intermediate[4095+3259:0+3259] + a; end
12'd3260: begin if(a[3260]==1) 
	 		intermediate[4095+3260:0+3260] <= intermediate[4095+3260:0+3260] + a; end
12'd3261: begin if(a[3261]==1) 
	 		intermediate[4095+3261:0+3261] <= intermediate[4095+3261:0+3261] + a; end
12'd3262: begin if(a[3262]==1) 
	 		intermediate[4095+3262:0+3262] <= intermediate[4095+3262:0+3262] + a; end
12'd3263: begin if(a[3263]==1) 
	 		intermediate[4095+3263:0+3263] <= intermediate[4095+3263:0+3263] + a; end
12'd3264: begin if(a[3264]==1) 
	 		intermediate[4095+3264:0+3264] <= intermediate[4095+3264:0+3264] + a; end
12'd3265: begin if(a[3265]==1) 
	 		intermediate[4095+3265:0+3265] <= intermediate[4095+3265:0+3265] + a; end
12'd3266: begin if(a[3266]==1) 
	 		intermediate[4095+3266:0+3266] <= intermediate[4095+3266:0+3266] + a; end
12'd3267: begin if(a[3267]==1) 
	 		intermediate[4095+3267:0+3267] <= intermediate[4095+3267:0+3267] + a; end
12'd3268: begin if(a[3268]==1) 
	 		intermediate[4095+3268:0+3268] <= intermediate[4095+3268:0+3268] + a; end
12'd3269: begin if(a[3269]==1) 
	 		intermediate[4095+3269:0+3269] <= intermediate[4095+3269:0+3269] + a; end
12'd3270: begin if(a[3270]==1) 
	 		intermediate[4095+3270:0+3270] <= intermediate[4095+3270:0+3270] + a; end
12'd3271: begin if(a[3271]==1) 
	 		intermediate[4095+3271:0+3271] <= intermediate[4095+3271:0+3271] + a; end
12'd3272: begin if(a[3272]==1) 
	 		intermediate[4095+3272:0+3272] <= intermediate[4095+3272:0+3272] + a; end
12'd3273: begin if(a[3273]==1) 
	 		intermediate[4095+3273:0+3273] <= intermediate[4095+3273:0+3273] + a; end
12'd3274: begin if(a[3274]==1) 
	 		intermediate[4095+3274:0+3274] <= intermediate[4095+3274:0+3274] + a; end
12'd3275: begin if(a[3275]==1) 
	 		intermediate[4095+3275:0+3275] <= intermediate[4095+3275:0+3275] + a; end
12'd3276: begin if(a[3276]==1) 
	 		intermediate[4095+3276:0+3276] <= intermediate[4095+3276:0+3276] + a; end
12'd3277: begin if(a[3277]==1) 
	 		intermediate[4095+3277:0+3277] <= intermediate[4095+3277:0+3277] + a; end
12'd3278: begin if(a[3278]==1) 
	 		intermediate[4095+3278:0+3278] <= intermediate[4095+3278:0+3278] + a; end
12'd3279: begin if(a[3279]==1) 
	 		intermediate[4095+3279:0+3279] <= intermediate[4095+3279:0+3279] + a; end
12'd3280: begin if(a[3280]==1) 
	 		intermediate[4095+3280:0+3280] <= intermediate[4095+3280:0+3280] + a; end
12'd3281: begin if(a[3281]==1) 
	 		intermediate[4095+3281:0+3281] <= intermediate[4095+3281:0+3281] + a; end
12'd3282: begin if(a[3282]==1) 
	 		intermediate[4095+3282:0+3282] <= intermediate[4095+3282:0+3282] + a; end
12'd3283: begin if(a[3283]==1) 
	 		intermediate[4095+3283:0+3283] <= intermediate[4095+3283:0+3283] + a; end
12'd3284: begin if(a[3284]==1) 
	 		intermediate[4095+3284:0+3284] <= intermediate[4095+3284:0+3284] + a; end
12'd3285: begin if(a[3285]==1) 
	 		intermediate[4095+3285:0+3285] <= intermediate[4095+3285:0+3285] + a; end
12'd3286: begin if(a[3286]==1) 
	 		intermediate[4095+3286:0+3286] <= intermediate[4095+3286:0+3286] + a; end
12'd3287: begin if(a[3287]==1) 
	 		intermediate[4095+3287:0+3287] <= intermediate[4095+3287:0+3287] + a; end
12'd3288: begin if(a[3288]==1) 
	 		intermediate[4095+3288:0+3288] <= intermediate[4095+3288:0+3288] + a; end
12'd3289: begin if(a[3289]==1) 
	 		intermediate[4095+3289:0+3289] <= intermediate[4095+3289:0+3289] + a; end
12'd3290: begin if(a[3290]==1) 
	 		intermediate[4095+3290:0+3290] <= intermediate[4095+3290:0+3290] + a; end
12'd3291: begin if(a[3291]==1) 
	 		intermediate[4095+3291:0+3291] <= intermediate[4095+3291:0+3291] + a; end
12'd3292: begin if(a[3292]==1) 
	 		intermediate[4095+3292:0+3292] <= intermediate[4095+3292:0+3292] + a; end
12'd3293: begin if(a[3293]==1) 
	 		intermediate[4095+3293:0+3293] <= intermediate[4095+3293:0+3293] + a; end
12'd3294: begin if(a[3294]==1) 
	 		intermediate[4095+3294:0+3294] <= intermediate[4095+3294:0+3294] + a; end
12'd3295: begin if(a[3295]==1) 
	 		intermediate[4095+3295:0+3295] <= intermediate[4095+3295:0+3295] + a; end
12'd3296: begin if(a[3296]==1) 
	 		intermediate[4095+3296:0+3296] <= intermediate[4095+3296:0+3296] + a; end
12'd3297: begin if(a[3297]==1) 
	 		intermediate[4095+3297:0+3297] <= intermediate[4095+3297:0+3297] + a; end
12'd3298: begin if(a[3298]==1) 
	 		intermediate[4095+3298:0+3298] <= intermediate[4095+3298:0+3298] + a; end
12'd3299: begin if(a[3299]==1) 
	 		intermediate[4095+3299:0+3299] <= intermediate[4095+3299:0+3299] + a; end
12'd3300: begin if(a[3300]==1) 
	 		intermediate[4095+3300:0+3300] <= intermediate[4095+3300:0+3300] + a; end
12'd3301: begin if(a[3301]==1) 
	 		intermediate[4095+3301:0+3301] <= intermediate[4095+3301:0+3301] + a; end
12'd3302: begin if(a[3302]==1) 
	 		intermediate[4095+3302:0+3302] <= intermediate[4095+3302:0+3302] + a; end
12'd3303: begin if(a[3303]==1) 
	 		intermediate[4095+3303:0+3303] <= intermediate[4095+3303:0+3303] + a; end
12'd3304: begin if(a[3304]==1) 
	 		intermediate[4095+3304:0+3304] <= intermediate[4095+3304:0+3304] + a; end
12'd3305: begin if(a[3305]==1) 
	 		intermediate[4095+3305:0+3305] <= intermediate[4095+3305:0+3305] + a; end
12'd3306: begin if(a[3306]==1) 
	 		intermediate[4095+3306:0+3306] <= intermediate[4095+3306:0+3306] + a; end
12'd3307: begin if(a[3307]==1) 
	 		intermediate[4095+3307:0+3307] <= intermediate[4095+3307:0+3307] + a; end
12'd3308: begin if(a[3308]==1) 
	 		intermediate[4095+3308:0+3308] <= intermediate[4095+3308:0+3308] + a; end
12'd3309: begin if(a[3309]==1) 
	 		intermediate[4095+3309:0+3309] <= intermediate[4095+3309:0+3309] + a; end
12'd3310: begin if(a[3310]==1) 
	 		intermediate[4095+3310:0+3310] <= intermediate[4095+3310:0+3310] + a; end
12'd3311: begin if(a[3311]==1) 
	 		intermediate[4095+3311:0+3311] <= intermediate[4095+3311:0+3311] + a; end
12'd3312: begin if(a[3312]==1) 
	 		intermediate[4095+3312:0+3312] <= intermediate[4095+3312:0+3312] + a; end
12'd3313: begin if(a[3313]==1) 
	 		intermediate[4095+3313:0+3313] <= intermediate[4095+3313:0+3313] + a; end
12'd3314: begin if(a[3314]==1) 
	 		intermediate[4095+3314:0+3314] <= intermediate[4095+3314:0+3314] + a; end
12'd3315: begin if(a[3315]==1) 
	 		intermediate[4095+3315:0+3315] <= intermediate[4095+3315:0+3315] + a; end
12'd3316: begin if(a[3316]==1) 
	 		intermediate[4095+3316:0+3316] <= intermediate[4095+3316:0+3316] + a; end
12'd3317: begin if(a[3317]==1) 
	 		intermediate[4095+3317:0+3317] <= intermediate[4095+3317:0+3317] + a; end
12'd3318: begin if(a[3318]==1) 
	 		intermediate[4095+3318:0+3318] <= intermediate[4095+3318:0+3318] + a; end
12'd3319: begin if(a[3319]==1) 
	 		intermediate[4095+3319:0+3319] <= intermediate[4095+3319:0+3319] + a; end
12'd3320: begin if(a[3320]==1) 
	 		intermediate[4095+3320:0+3320] <= intermediate[4095+3320:0+3320] + a; end
12'd3321: begin if(a[3321]==1) 
	 		intermediate[4095+3321:0+3321] <= intermediate[4095+3321:0+3321] + a; end
12'd3322: begin if(a[3322]==1) 
	 		intermediate[4095+3322:0+3322] <= intermediate[4095+3322:0+3322] + a; end
12'd3323: begin if(a[3323]==1) 
	 		intermediate[4095+3323:0+3323] <= intermediate[4095+3323:0+3323] + a; end
12'd3324: begin if(a[3324]==1) 
	 		intermediate[4095+3324:0+3324] <= intermediate[4095+3324:0+3324] + a; end
12'd3325: begin if(a[3325]==1) 
	 		intermediate[4095+3325:0+3325] <= intermediate[4095+3325:0+3325] + a; end
12'd3326: begin if(a[3326]==1) 
	 		intermediate[4095+3326:0+3326] <= intermediate[4095+3326:0+3326] + a; end
12'd3327: begin if(a[3327]==1) 
	 		intermediate[4095+3327:0+3327] <= intermediate[4095+3327:0+3327] + a; end
12'd3328: begin if(a[3328]==1) 
	 		intermediate[4095+3328:0+3328] <= intermediate[4095+3328:0+3328] + a; end
12'd3329: begin if(a[3329]==1) 
	 		intermediate[4095+3329:0+3329] <= intermediate[4095+3329:0+3329] + a; end
12'd3330: begin if(a[3330]==1) 
	 		intermediate[4095+3330:0+3330] <= intermediate[4095+3330:0+3330] + a; end
12'd3331: begin if(a[3331]==1) 
	 		intermediate[4095+3331:0+3331] <= intermediate[4095+3331:0+3331] + a; end
12'd3332: begin if(a[3332]==1) 
	 		intermediate[4095+3332:0+3332] <= intermediate[4095+3332:0+3332] + a; end
12'd3333: begin if(a[3333]==1) 
	 		intermediate[4095+3333:0+3333] <= intermediate[4095+3333:0+3333] + a; end
12'd3334: begin if(a[3334]==1) 
	 		intermediate[4095+3334:0+3334] <= intermediate[4095+3334:0+3334] + a; end
12'd3335: begin if(a[3335]==1) 
	 		intermediate[4095+3335:0+3335] <= intermediate[4095+3335:0+3335] + a; end
12'd3336: begin if(a[3336]==1) 
	 		intermediate[4095+3336:0+3336] <= intermediate[4095+3336:0+3336] + a; end
12'd3337: begin if(a[3337]==1) 
	 		intermediate[4095+3337:0+3337] <= intermediate[4095+3337:0+3337] + a; end
12'd3338: begin if(a[3338]==1) 
	 		intermediate[4095+3338:0+3338] <= intermediate[4095+3338:0+3338] + a; end
12'd3339: begin if(a[3339]==1) 
	 		intermediate[4095+3339:0+3339] <= intermediate[4095+3339:0+3339] + a; end
12'd3340: begin if(a[3340]==1) 
	 		intermediate[4095+3340:0+3340] <= intermediate[4095+3340:0+3340] + a; end
12'd3341: begin if(a[3341]==1) 
	 		intermediate[4095+3341:0+3341] <= intermediate[4095+3341:0+3341] + a; end
12'd3342: begin if(a[3342]==1) 
	 		intermediate[4095+3342:0+3342] <= intermediate[4095+3342:0+3342] + a; end
12'd3343: begin if(a[3343]==1) 
	 		intermediate[4095+3343:0+3343] <= intermediate[4095+3343:0+3343] + a; end
12'd3344: begin if(a[3344]==1) 
	 		intermediate[4095+3344:0+3344] <= intermediate[4095+3344:0+3344] + a; end
12'd3345: begin if(a[3345]==1) 
	 		intermediate[4095+3345:0+3345] <= intermediate[4095+3345:0+3345] + a; end
12'd3346: begin if(a[3346]==1) 
	 		intermediate[4095+3346:0+3346] <= intermediate[4095+3346:0+3346] + a; end
12'd3347: begin if(a[3347]==1) 
	 		intermediate[4095+3347:0+3347] <= intermediate[4095+3347:0+3347] + a; end
12'd3348: begin if(a[3348]==1) 
	 		intermediate[4095+3348:0+3348] <= intermediate[4095+3348:0+3348] + a; end
12'd3349: begin if(a[3349]==1) 
	 		intermediate[4095+3349:0+3349] <= intermediate[4095+3349:0+3349] + a; end
12'd3350: begin if(a[3350]==1) 
	 		intermediate[4095+3350:0+3350] <= intermediate[4095+3350:0+3350] + a; end
12'd3351: begin if(a[3351]==1) 
	 		intermediate[4095+3351:0+3351] <= intermediate[4095+3351:0+3351] + a; end
12'd3352: begin if(a[3352]==1) 
	 		intermediate[4095+3352:0+3352] <= intermediate[4095+3352:0+3352] + a; end
12'd3353: begin if(a[3353]==1) 
	 		intermediate[4095+3353:0+3353] <= intermediate[4095+3353:0+3353] + a; end
12'd3354: begin if(a[3354]==1) 
	 		intermediate[4095+3354:0+3354] <= intermediate[4095+3354:0+3354] + a; end
12'd3355: begin if(a[3355]==1) 
	 		intermediate[4095+3355:0+3355] <= intermediate[4095+3355:0+3355] + a; end
12'd3356: begin if(a[3356]==1) 
	 		intermediate[4095+3356:0+3356] <= intermediate[4095+3356:0+3356] + a; end
12'd3357: begin if(a[3357]==1) 
	 		intermediate[4095+3357:0+3357] <= intermediate[4095+3357:0+3357] + a; end
12'd3358: begin if(a[3358]==1) 
	 		intermediate[4095+3358:0+3358] <= intermediate[4095+3358:0+3358] + a; end
12'd3359: begin if(a[3359]==1) 
	 		intermediate[4095+3359:0+3359] <= intermediate[4095+3359:0+3359] + a; end
12'd3360: begin if(a[3360]==1) 
	 		intermediate[4095+3360:0+3360] <= intermediate[4095+3360:0+3360] + a; end
12'd3361: begin if(a[3361]==1) 
	 		intermediate[4095+3361:0+3361] <= intermediate[4095+3361:0+3361] + a; end
12'd3362: begin if(a[3362]==1) 
	 		intermediate[4095+3362:0+3362] <= intermediate[4095+3362:0+3362] + a; end
12'd3363: begin if(a[3363]==1) 
	 		intermediate[4095+3363:0+3363] <= intermediate[4095+3363:0+3363] + a; end
12'd3364: begin if(a[3364]==1) 
	 		intermediate[4095+3364:0+3364] <= intermediate[4095+3364:0+3364] + a; end
12'd3365: begin if(a[3365]==1) 
	 		intermediate[4095+3365:0+3365] <= intermediate[4095+3365:0+3365] + a; end
12'd3366: begin if(a[3366]==1) 
	 		intermediate[4095+3366:0+3366] <= intermediate[4095+3366:0+3366] + a; end
12'd3367: begin if(a[3367]==1) 
	 		intermediate[4095+3367:0+3367] <= intermediate[4095+3367:0+3367] + a; end
12'd3368: begin if(a[3368]==1) 
	 		intermediate[4095+3368:0+3368] <= intermediate[4095+3368:0+3368] + a; end
12'd3369: begin if(a[3369]==1) 
	 		intermediate[4095+3369:0+3369] <= intermediate[4095+3369:0+3369] + a; end
12'd3370: begin if(a[3370]==1) 
	 		intermediate[4095+3370:0+3370] <= intermediate[4095+3370:0+3370] + a; end
12'd3371: begin if(a[3371]==1) 
	 		intermediate[4095+3371:0+3371] <= intermediate[4095+3371:0+3371] + a; end
12'd3372: begin if(a[3372]==1) 
	 		intermediate[4095+3372:0+3372] <= intermediate[4095+3372:0+3372] + a; end
12'd3373: begin if(a[3373]==1) 
	 		intermediate[4095+3373:0+3373] <= intermediate[4095+3373:0+3373] + a; end
12'd3374: begin if(a[3374]==1) 
	 		intermediate[4095+3374:0+3374] <= intermediate[4095+3374:0+3374] + a; end
12'd3375: begin if(a[3375]==1) 
	 		intermediate[4095+3375:0+3375] <= intermediate[4095+3375:0+3375] + a; end
12'd3376: begin if(a[3376]==1) 
	 		intermediate[4095+3376:0+3376] <= intermediate[4095+3376:0+3376] + a; end
12'd3377: begin if(a[3377]==1) 
	 		intermediate[4095+3377:0+3377] <= intermediate[4095+3377:0+3377] + a; end
12'd3378: begin if(a[3378]==1) 
	 		intermediate[4095+3378:0+3378] <= intermediate[4095+3378:0+3378] + a; end
12'd3379: begin if(a[3379]==1) 
	 		intermediate[4095+3379:0+3379] <= intermediate[4095+3379:0+3379] + a; end
12'd3380: begin if(a[3380]==1) 
	 		intermediate[4095+3380:0+3380] <= intermediate[4095+3380:0+3380] + a; end
12'd3381: begin if(a[3381]==1) 
	 		intermediate[4095+3381:0+3381] <= intermediate[4095+3381:0+3381] + a; end
12'd3382: begin if(a[3382]==1) 
	 		intermediate[4095+3382:0+3382] <= intermediate[4095+3382:0+3382] + a; end
12'd3383: begin if(a[3383]==1) 
	 		intermediate[4095+3383:0+3383] <= intermediate[4095+3383:0+3383] + a; end
12'd3384: begin if(a[3384]==1) 
	 		intermediate[4095+3384:0+3384] <= intermediate[4095+3384:0+3384] + a; end
12'd3385: begin if(a[3385]==1) 
	 		intermediate[4095+3385:0+3385] <= intermediate[4095+3385:0+3385] + a; end
12'd3386: begin if(a[3386]==1) 
	 		intermediate[4095+3386:0+3386] <= intermediate[4095+3386:0+3386] + a; end
12'd3387: begin if(a[3387]==1) 
	 		intermediate[4095+3387:0+3387] <= intermediate[4095+3387:0+3387] + a; end
12'd3388: begin if(a[3388]==1) 
	 		intermediate[4095+3388:0+3388] <= intermediate[4095+3388:0+3388] + a; end
12'd3389: begin if(a[3389]==1) 
	 		intermediate[4095+3389:0+3389] <= intermediate[4095+3389:0+3389] + a; end
12'd3390: begin if(a[3390]==1) 
	 		intermediate[4095+3390:0+3390] <= intermediate[4095+3390:0+3390] + a; end
12'd3391: begin if(a[3391]==1) 
	 		intermediate[4095+3391:0+3391] <= intermediate[4095+3391:0+3391] + a; end
12'd3392: begin if(a[3392]==1) 
	 		intermediate[4095+3392:0+3392] <= intermediate[4095+3392:0+3392] + a; end
12'd3393: begin if(a[3393]==1) 
	 		intermediate[4095+3393:0+3393] <= intermediate[4095+3393:0+3393] + a; end
12'd3394: begin if(a[3394]==1) 
	 		intermediate[4095+3394:0+3394] <= intermediate[4095+3394:0+3394] + a; end
12'd3395: begin if(a[3395]==1) 
	 		intermediate[4095+3395:0+3395] <= intermediate[4095+3395:0+3395] + a; end
12'd3396: begin if(a[3396]==1) 
	 		intermediate[4095+3396:0+3396] <= intermediate[4095+3396:0+3396] + a; end
12'd3397: begin if(a[3397]==1) 
	 		intermediate[4095+3397:0+3397] <= intermediate[4095+3397:0+3397] + a; end
12'd3398: begin if(a[3398]==1) 
	 		intermediate[4095+3398:0+3398] <= intermediate[4095+3398:0+3398] + a; end
12'd3399: begin if(a[3399]==1) 
	 		intermediate[4095+3399:0+3399] <= intermediate[4095+3399:0+3399] + a; end
12'd3400: begin if(a[3400]==1) 
	 		intermediate[4095+3400:0+3400] <= intermediate[4095+3400:0+3400] + a; end
12'd3401: begin if(a[3401]==1) 
	 		intermediate[4095+3401:0+3401] <= intermediate[4095+3401:0+3401] + a; end
12'd3402: begin if(a[3402]==1) 
	 		intermediate[4095+3402:0+3402] <= intermediate[4095+3402:0+3402] + a; end
12'd3403: begin if(a[3403]==1) 
	 		intermediate[4095+3403:0+3403] <= intermediate[4095+3403:0+3403] + a; end
12'd3404: begin if(a[3404]==1) 
	 		intermediate[4095+3404:0+3404] <= intermediate[4095+3404:0+3404] + a; end
12'd3405: begin if(a[3405]==1) 
	 		intermediate[4095+3405:0+3405] <= intermediate[4095+3405:0+3405] + a; end
12'd3406: begin if(a[3406]==1) 
	 		intermediate[4095+3406:0+3406] <= intermediate[4095+3406:0+3406] + a; end
12'd3407: begin if(a[3407]==1) 
	 		intermediate[4095+3407:0+3407] <= intermediate[4095+3407:0+3407] + a; end
12'd3408: begin if(a[3408]==1) 
	 		intermediate[4095+3408:0+3408] <= intermediate[4095+3408:0+3408] + a; end
12'd3409: begin if(a[3409]==1) 
	 		intermediate[4095+3409:0+3409] <= intermediate[4095+3409:0+3409] + a; end
12'd3410: begin if(a[3410]==1) 
	 		intermediate[4095+3410:0+3410] <= intermediate[4095+3410:0+3410] + a; end
12'd3411: begin if(a[3411]==1) 
	 		intermediate[4095+3411:0+3411] <= intermediate[4095+3411:0+3411] + a; end
12'd3412: begin if(a[3412]==1) 
	 		intermediate[4095+3412:0+3412] <= intermediate[4095+3412:0+3412] + a; end
12'd3413: begin if(a[3413]==1) 
	 		intermediate[4095+3413:0+3413] <= intermediate[4095+3413:0+3413] + a; end
12'd3414: begin if(a[3414]==1) 
	 		intermediate[4095+3414:0+3414] <= intermediate[4095+3414:0+3414] + a; end
12'd3415: begin if(a[3415]==1) 
	 		intermediate[4095+3415:0+3415] <= intermediate[4095+3415:0+3415] + a; end
12'd3416: begin if(a[3416]==1) 
	 		intermediate[4095+3416:0+3416] <= intermediate[4095+3416:0+3416] + a; end
12'd3417: begin if(a[3417]==1) 
	 		intermediate[4095+3417:0+3417] <= intermediate[4095+3417:0+3417] + a; end
12'd3418: begin if(a[3418]==1) 
	 		intermediate[4095+3418:0+3418] <= intermediate[4095+3418:0+3418] + a; end
12'd3419: begin if(a[3419]==1) 
	 		intermediate[4095+3419:0+3419] <= intermediate[4095+3419:0+3419] + a; end
12'd3420: begin if(a[3420]==1) 
	 		intermediate[4095+3420:0+3420] <= intermediate[4095+3420:0+3420] + a; end
12'd3421: begin if(a[3421]==1) 
	 		intermediate[4095+3421:0+3421] <= intermediate[4095+3421:0+3421] + a; end
12'd3422: begin if(a[3422]==1) 
	 		intermediate[4095+3422:0+3422] <= intermediate[4095+3422:0+3422] + a; end
12'd3423: begin if(a[3423]==1) 
	 		intermediate[4095+3423:0+3423] <= intermediate[4095+3423:0+3423] + a; end
12'd3424: begin if(a[3424]==1) 
	 		intermediate[4095+3424:0+3424] <= intermediate[4095+3424:0+3424] + a; end
12'd3425: begin if(a[3425]==1) 
	 		intermediate[4095+3425:0+3425] <= intermediate[4095+3425:0+3425] + a; end
12'd3426: begin if(a[3426]==1) 
	 		intermediate[4095+3426:0+3426] <= intermediate[4095+3426:0+3426] + a; end
12'd3427: begin if(a[3427]==1) 
	 		intermediate[4095+3427:0+3427] <= intermediate[4095+3427:0+3427] + a; end
12'd3428: begin if(a[3428]==1) 
	 		intermediate[4095+3428:0+3428] <= intermediate[4095+3428:0+3428] + a; end
12'd3429: begin if(a[3429]==1) 
	 		intermediate[4095+3429:0+3429] <= intermediate[4095+3429:0+3429] + a; end
12'd3430: begin if(a[3430]==1) 
	 		intermediate[4095+3430:0+3430] <= intermediate[4095+3430:0+3430] + a; end
12'd3431: begin if(a[3431]==1) 
	 		intermediate[4095+3431:0+3431] <= intermediate[4095+3431:0+3431] + a; end
12'd3432: begin if(a[3432]==1) 
	 		intermediate[4095+3432:0+3432] <= intermediate[4095+3432:0+3432] + a; end
12'd3433: begin if(a[3433]==1) 
	 		intermediate[4095+3433:0+3433] <= intermediate[4095+3433:0+3433] + a; end
12'd3434: begin if(a[3434]==1) 
	 		intermediate[4095+3434:0+3434] <= intermediate[4095+3434:0+3434] + a; end
12'd3435: begin if(a[3435]==1) 
	 		intermediate[4095+3435:0+3435] <= intermediate[4095+3435:0+3435] + a; end
12'd3436: begin if(a[3436]==1) 
	 		intermediate[4095+3436:0+3436] <= intermediate[4095+3436:0+3436] + a; end
12'd3437: begin if(a[3437]==1) 
	 		intermediate[4095+3437:0+3437] <= intermediate[4095+3437:0+3437] + a; end
12'd3438: begin if(a[3438]==1) 
	 		intermediate[4095+3438:0+3438] <= intermediate[4095+3438:0+3438] + a; end
12'd3439: begin if(a[3439]==1) 
	 		intermediate[4095+3439:0+3439] <= intermediate[4095+3439:0+3439] + a; end
12'd3440: begin if(a[3440]==1) 
	 		intermediate[4095+3440:0+3440] <= intermediate[4095+3440:0+3440] + a; end
12'd3441: begin if(a[3441]==1) 
	 		intermediate[4095+3441:0+3441] <= intermediate[4095+3441:0+3441] + a; end
12'd3442: begin if(a[3442]==1) 
	 		intermediate[4095+3442:0+3442] <= intermediate[4095+3442:0+3442] + a; end
12'd3443: begin if(a[3443]==1) 
	 		intermediate[4095+3443:0+3443] <= intermediate[4095+3443:0+3443] + a; end
12'd3444: begin if(a[3444]==1) 
	 		intermediate[4095+3444:0+3444] <= intermediate[4095+3444:0+3444] + a; end
12'd3445: begin if(a[3445]==1) 
	 		intermediate[4095+3445:0+3445] <= intermediate[4095+3445:0+3445] + a; end
12'd3446: begin if(a[3446]==1) 
	 		intermediate[4095+3446:0+3446] <= intermediate[4095+3446:0+3446] + a; end
12'd3447: begin if(a[3447]==1) 
	 		intermediate[4095+3447:0+3447] <= intermediate[4095+3447:0+3447] + a; end
12'd3448: begin if(a[3448]==1) 
	 		intermediate[4095+3448:0+3448] <= intermediate[4095+3448:0+3448] + a; end
12'd3449: begin if(a[3449]==1) 
	 		intermediate[4095+3449:0+3449] <= intermediate[4095+3449:0+3449] + a; end
12'd3450: begin if(a[3450]==1) 
	 		intermediate[4095+3450:0+3450] <= intermediate[4095+3450:0+3450] + a; end
12'd3451: begin if(a[3451]==1) 
	 		intermediate[4095+3451:0+3451] <= intermediate[4095+3451:0+3451] + a; end
12'd3452: begin if(a[3452]==1) 
	 		intermediate[4095+3452:0+3452] <= intermediate[4095+3452:0+3452] + a; end
12'd3453: begin if(a[3453]==1) 
	 		intermediate[4095+3453:0+3453] <= intermediate[4095+3453:0+3453] + a; end
12'd3454: begin if(a[3454]==1) 
	 		intermediate[4095+3454:0+3454] <= intermediate[4095+3454:0+3454] + a; end
12'd3455: begin if(a[3455]==1) 
	 		intermediate[4095+3455:0+3455] <= intermediate[4095+3455:0+3455] + a; end
12'd3456: begin if(a[3456]==1) 
	 		intermediate[4095+3456:0+3456] <= intermediate[4095+3456:0+3456] + a; end
12'd3457: begin if(a[3457]==1) 
	 		intermediate[4095+3457:0+3457] <= intermediate[4095+3457:0+3457] + a; end
12'd3458: begin if(a[3458]==1) 
	 		intermediate[4095+3458:0+3458] <= intermediate[4095+3458:0+3458] + a; end
12'd3459: begin if(a[3459]==1) 
	 		intermediate[4095+3459:0+3459] <= intermediate[4095+3459:0+3459] + a; end
12'd3460: begin if(a[3460]==1) 
	 		intermediate[4095+3460:0+3460] <= intermediate[4095+3460:0+3460] + a; end
12'd3461: begin if(a[3461]==1) 
	 		intermediate[4095+3461:0+3461] <= intermediate[4095+3461:0+3461] + a; end
12'd3462: begin if(a[3462]==1) 
	 		intermediate[4095+3462:0+3462] <= intermediate[4095+3462:0+3462] + a; end
12'd3463: begin if(a[3463]==1) 
	 		intermediate[4095+3463:0+3463] <= intermediate[4095+3463:0+3463] + a; end
12'd3464: begin if(a[3464]==1) 
	 		intermediate[4095+3464:0+3464] <= intermediate[4095+3464:0+3464] + a; end
12'd3465: begin if(a[3465]==1) 
	 		intermediate[4095+3465:0+3465] <= intermediate[4095+3465:0+3465] + a; end
12'd3466: begin if(a[3466]==1) 
	 		intermediate[4095+3466:0+3466] <= intermediate[4095+3466:0+3466] + a; end
12'd3467: begin if(a[3467]==1) 
	 		intermediate[4095+3467:0+3467] <= intermediate[4095+3467:0+3467] + a; end
12'd3468: begin if(a[3468]==1) 
	 		intermediate[4095+3468:0+3468] <= intermediate[4095+3468:0+3468] + a; end
12'd3469: begin if(a[3469]==1) 
	 		intermediate[4095+3469:0+3469] <= intermediate[4095+3469:0+3469] + a; end
12'd3470: begin if(a[3470]==1) 
	 		intermediate[4095+3470:0+3470] <= intermediate[4095+3470:0+3470] + a; end
12'd3471: begin if(a[3471]==1) 
	 		intermediate[4095+3471:0+3471] <= intermediate[4095+3471:0+3471] + a; end
12'd3472: begin if(a[3472]==1) 
	 		intermediate[4095+3472:0+3472] <= intermediate[4095+3472:0+3472] + a; end
12'd3473: begin if(a[3473]==1) 
	 		intermediate[4095+3473:0+3473] <= intermediate[4095+3473:0+3473] + a; end
12'd3474: begin if(a[3474]==1) 
	 		intermediate[4095+3474:0+3474] <= intermediate[4095+3474:0+3474] + a; end
12'd3475: begin if(a[3475]==1) 
	 		intermediate[4095+3475:0+3475] <= intermediate[4095+3475:0+3475] + a; end
12'd3476: begin if(a[3476]==1) 
	 		intermediate[4095+3476:0+3476] <= intermediate[4095+3476:0+3476] + a; end
12'd3477: begin if(a[3477]==1) 
	 		intermediate[4095+3477:0+3477] <= intermediate[4095+3477:0+3477] + a; end
12'd3478: begin if(a[3478]==1) 
	 		intermediate[4095+3478:0+3478] <= intermediate[4095+3478:0+3478] + a; end
12'd3479: begin if(a[3479]==1) 
	 		intermediate[4095+3479:0+3479] <= intermediate[4095+3479:0+3479] + a; end
12'd3480: begin if(a[3480]==1) 
	 		intermediate[4095+3480:0+3480] <= intermediate[4095+3480:0+3480] + a; end
12'd3481: begin if(a[3481]==1) 
	 		intermediate[4095+3481:0+3481] <= intermediate[4095+3481:0+3481] + a; end
12'd3482: begin if(a[3482]==1) 
	 		intermediate[4095+3482:0+3482] <= intermediate[4095+3482:0+3482] + a; end
12'd3483: begin if(a[3483]==1) 
	 		intermediate[4095+3483:0+3483] <= intermediate[4095+3483:0+3483] + a; end
12'd3484: begin if(a[3484]==1) 
	 		intermediate[4095+3484:0+3484] <= intermediate[4095+3484:0+3484] + a; end
12'd3485: begin if(a[3485]==1) 
	 		intermediate[4095+3485:0+3485] <= intermediate[4095+3485:0+3485] + a; end
12'd3486: begin if(a[3486]==1) 
	 		intermediate[4095+3486:0+3486] <= intermediate[4095+3486:0+3486] + a; end
12'd3487: begin if(a[3487]==1) 
	 		intermediate[4095+3487:0+3487] <= intermediate[4095+3487:0+3487] + a; end
12'd3488: begin if(a[3488]==1) 
	 		intermediate[4095+3488:0+3488] <= intermediate[4095+3488:0+3488] + a; end
12'd3489: begin if(a[3489]==1) 
	 		intermediate[4095+3489:0+3489] <= intermediate[4095+3489:0+3489] + a; end
12'd3490: begin if(a[3490]==1) 
	 		intermediate[4095+3490:0+3490] <= intermediate[4095+3490:0+3490] + a; end
12'd3491: begin if(a[3491]==1) 
	 		intermediate[4095+3491:0+3491] <= intermediate[4095+3491:0+3491] + a; end
12'd3492: begin if(a[3492]==1) 
	 		intermediate[4095+3492:0+3492] <= intermediate[4095+3492:0+3492] + a; end
12'd3493: begin if(a[3493]==1) 
	 		intermediate[4095+3493:0+3493] <= intermediate[4095+3493:0+3493] + a; end
12'd3494: begin if(a[3494]==1) 
	 		intermediate[4095+3494:0+3494] <= intermediate[4095+3494:0+3494] + a; end
12'd3495: begin if(a[3495]==1) 
	 		intermediate[4095+3495:0+3495] <= intermediate[4095+3495:0+3495] + a; end
12'd3496: begin if(a[3496]==1) 
	 		intermediate[4095+3496:0+3496] <= intermediate[4095+3496:0+3496] + a; end
12'd3497: begin if(a[3497]==1) 
	 		intermediate[4095+3497:0+3497] <= intermediate[4095+3497:0+3497] + a; end
12'd3498: begin if(a[3498]==1) 
	 		intermediate[4095+3498:0+3498] <= intermediate[4095+3498:0+3498] + a; end
12'd3499: begin if(a[3499]==1) 
	 		intermediate[4095+3499:0+3499] <= intermediate[4095+3499:0+3499] + a; end
12'd3500: begin if(a[3500]==1) 
	 		intermediate[4095+3500:0+3500] <= intermediate[4095+3500:0+3500] + a; end
12'd3501: begin if(a[3501]==1) 
	 		intermediate[4095+3501:0+3501] <= intermediate[4095+3501:0+3501] + a; end
12'd3502: begin if(a[3502]==1) 
	 		intermediate[4095+3502:0+3502] <= intermediate[4095+3502:0+3502] + a; end
12'd3503: begin if(a[3503]==1) 
	 		intermediate[4095+3503:0+3503] <= intermediate[4095+3503:0+3503] + a; end
12'd3504: begin if(a[3504]==1) 
	 		intermediate[4095+3504:0+3504] <= intermediate[4095+3504:0+3504] + a; end
12'd3505: begin if(a[3505]==1) 
	 		intermediate[4095+3505:0+3505] <= intermediate[4095+3505:0+3505] + a; end
12'd3506: begin if(a[3506]==1) 
	 		intermediate[4095+3506:0+3506] <= intermediate[4095+3506:0+3506] + a; end
12'd3507: begin if(a[3507]==1) 
	 		intermediate[4095+3507:0+3507] <= intermediate[4095+3507:0+3507] + a; end
12'd3508: begin if(a[3508]==1) 
	 		intermediate[4095+3508:0+3508] <= intermediate[4095+3508:0+3508] + a; end
12'd3509: begin if(a[3509]==1) 
	 		intermediate[4095+3509:0+3509] <= intermediate[4095+3509:0+3509] + a; end
12'd3510: begin if(a[3510]==1) 
	 		intermediate[4095+3510:0+3510] <= intermediate[4095+3510:0+3510] + a; end
12'd3511: begin if(a[3511]==1) 
	 		intermediate[4095+3511:0+3511] <= intermediate[4095+3511:0+3511] + a; end
12'd3512: begin if(a[3512]==1) 
	 		intermediate[4095+3512:0+3512] <= intermediate[4095+3512:0+3512] + a; end
12'd3513: begin if(a[3513]==1) 
	 		intermediate[4095+3513:0+3513] <= intermediate[4095+3513:0+3513] + a; end
12'd3514: begin if(a[3514]==1) 
	 		intermediate[4095+3514:0+3514] <= intermediate[4095+3514:0+3514] + a; end
12'd3515: begin if(a[3515]==1) 
	 		intermediate[4095+3515:0+3515] <= intermediate[4095+3515:0+3515] + a; end
12'd3516: begin if(a[3516]==1) 
	 		intermediate[4095+3516:0+3516] <= intermediate[4095+3516:0+3516] + a; end
12'd3517: begin if(a[3517]==1) 
	 		intermediate[4095+3517:0+3517] <= intermediate[4095+3517:0+3517] + a; end
12'd3518: begin if(a[3518]==1) 
	 		intermediate[4095+3518:0+3518] <= intermediate[4095+3518:0+3518] + a; end
12'd3519: begin if(a[3519]==1) 
	 		intermediate[4095+3519:0+3519] <= intermediate[4095+3519:0+3519] + a; end
12'd3520: begin if(a[3520]==1) 
	 		intermediate[4095+3520:0+3520] <= intermediate[4095+3520:0+3520] + a; end
12'd3521: begin if(a[3521]==1) 
	 		intermediate[4095+3521:0+3521] <= intermediate[4095+3521:0+3521] + a; end
12'd3522: begin if(a[3522]==1) 
	 		intermediate[4095+3522:0+3522] <= intermediate[4095+3522:0+3522] + a; end
12'd3523: begin if(a[3523]==1) 
	 		intermediate[4095+3523:0+3523] <= intermediate[4095+3523:0+3523] + a; end
12'd3524: begin if(a[3524]==1) 
	 		intermediate[4095+3524:0+3524] <= intermediate[4095+3524:0+3524] + a; end
12'd3525: begin if(a[3525]==1) 
	 		intermediate[4095+3525:0+3525] <= intermediate[4095+3525:0+3525] + a; end
12'd3526: begin if(a[3526]==1) 
	 		intermediate[4095+3526:0+3526] <= intermediate[4095+3526:0+3526] + a; end
12'd3527: begin if(a[3527]==1) 
	 		intermediate[4095+3527:0+3527] <= intermediate[4095+3527:0+3527] + a; end
12'd3528: begin if(a[3528]==1) 
	 		intermediate[4095+3528:0+3528] <= intermediate[4095+3528:0+3528] + a; end
12'd3529: begin if(a[3529]==1) 
	 		intermediate[4095+3529:0+3529] <= intermediate[4095+3529:0+3529] + a; end
12'd3530: begin if(a[3530]==1) 
	 		intermediate[4095+3530:0+3530] <= intermediate[4095+3530:0+3530] + a; end
12'd3531: begin if(a[3531]==1) 
	 		intermediate[4095+3531:0+3531] <= intermediate[4095+3531:0+3531] + a; end
12'd3532: begin if(a[3532]==1) 
	 		intermediate[4095+3532:0+3532] <= intermediate[4095+3532:0+3532] + a; end
12'd3533: begin if(a[3533]==1) 
	 		intermediate[4095+3533:0+3533] <= intermediate[4095+3533:0+3533] + a; end
12'd3534: begin if(a[3534]==1) 
	 		intermediate[4095+3534:0+3534] <= intermediate[4095+3534:0+3534] + a; end
12'd3535: begin if(a[3535]==1) 
	 		intermediate[4095+3535:0+3535] <= intermediate[4095+3535:0+3535] + a; end
12'd3536: begin if(a[3536]==1) 
	 		intermediate[4095+3536:0+3536] <= intermediate[4095+3536:0+3536] + a; end
12'd3537: begin if(a[3537]==1) 
	 		intermediate[4095+3537:0+3537] <= intermediate[4095+3537:0+3537] + a; end
12'd3538: begin if(a[3538]==1) 
	 		intermediate[4095+3538:0+3538] <= intermediate[4095+3538:0+3538] + a; end
12'd3539: begin if(a[3539]==1) 
	 		intermediate[4095+3539:0+3539] <= intermediate[4095+3539:0+3539] + a; end
12'd3540: begin if(a[3540]==1) 
	 		intermediate[4095+3540:0+3540] <= intermediate[4095+3540:0+3540] + a; end
12'd3541: begin if(a[3541]==1) 
	 		intermediate[4095+3541:0+3541] <= intermediate[4095+3541:0+3541] + a; end
12'd3542: begin if(a[3542]==1) 
	 		intermediate[4095+3542:0+3542] <= intermediate[4095+3542:0+3542] + a; end
12'd3543: begin if(a[3543]==1) 
	 		intermediate[4095+3543:0+3543] <= intermediate[4095+3543:0+3543] + a; end
12'd3544: begin if(a[3544]==1) 
	 		intermediate[4095+3544:0+3544] <= intermediate[4095+3544:0+3544] + a; end
12'd3545: begin if(a[3545]==1) 
	 		intermediate[4095+3545:0+3545] <= intermediate[4095+3545:0+3545] + a; end
12'd3546: begin if(a[3546]==1) 
	 		intermediate[4095+3546:0+3546] <= intermediate[4095+3546:0+3546] + a; end
12'd3547: begin if(a[3547]==1) 
	 		intermediate[4095+3547:0+3547] <= intermediate[4095+3547:0+3547] + a; end
12'd3548: begin if(a[3548]==1) 
	 		intermediate[4095+3548:0+3548] <= intermediate[4095+3548:0+3548] + a; end
12'd3549: begin if(a[3549]==1) 
	 		intermediate[4095+3549:0+3549] <= intermediate[4095+3549:0+3549] + a; end
12'd3550: begin if(a[3550]==1) 
	 		intermediate[4095+3550:0+3550] <= intermediate[4095+3550:0+3550] + a; end
12'd3551: begin if(a[3551]==1) 
	 		intermediate[4095+3551:0+3551] <= intermediate[4095+3551:0+3551] + a; end
12'd3552: begin if(a[3552]==1) 
	 		intermediate[4095+3552:0+3552] <= intermediate[4095+3552:0+3552] + a; end
12'd3553: begin if(a[3553]==1) 
	 		intermediate[4095+3553:0+3553] <= intermediate[4095+3553:0+3553] + a; end
12'd3554: begin if(a[3554]==1) 
	 		intermediate[4095+3554:0+3554] <= intermediate[4095+3554:0+3554] + a; end
12'd3555: begin if(a[3555]==1) 
	 		intermediate[4095+3555:0+3555] <= intermediate[4095+3555:0+3555] + a; end
12'd3556: begin if(a[3556]==1) 
	 		intermediate[4095+3556:0+3556] <= intermediate[4095+3556:0+3556] + a; end
12'd3557: begin if(a[3557]==1) 
	 		intermediate[4095+3557:0+3557] <= intermediate[4095+3557:0+3557] + a; end
12'd3558: begin if(a[3558]==1) 
	 		intermediate[4095+3558:0+3558] <= intermediate[4095+3558:0+3558] + a; end
12'd3559: begin if(a[3559]==1) 
	 		intermediate[4095+3559:0+3559] <= intermediate[4095+3559:0+3559] + a; end
12'd3560: begin if(a[3560]==1) 
	 		intermediate[4095+3560:0+3560] <= intermediate[4095+3560:0+3560] + a; end
12'd3561: begin if(a[3561]==1) 
	 		intermediate[4095+3561:0+3561] <= intermediate[4095+3561:0+3561] + a; end
12'd3562: begin if(a[3562]==1) 
	 		intermediate[4095+3562:0+3562] <= intermediate[4095+3562:0+3562] + a; end
12'd3563: begin if(a[3563]==1) 
	 		intermediate[4095+3563:0+3563] <= intermediate[4095+3563:0+3563] + a; end
12'd3564: begin if(a[3564]==1) 
	 		intermediate[4095+3564:0+3564] <= intermediate[4095+3564:0+3564] + a; end
12'd3565: begin if(a[3565]==1) 
	 		intermediate[4095+3565:0+3565] <= intermediate[4095+3565:0+3565] + a; end
12'd3566: begin if(a[3566]==1) 
	 		intermediate[4095+3566:0+3566] <= intermediate[4095+3566:0+3566] + a; end
12'd3567: begin if(a[3567]==1) 
	 		intermediate[4095+3567:0+3567] <= intermediate[4095+3567:0+3567] + a; end
12'd3568: begin if(a[3568]==1) 
	 		intermediate[4095+3568:0+3568] <= intermediate[4095+3568:0+3568] + a; end
12'd3569: begin if(a[3569]==1) 
	 		intermediate[4095+3569:0+3569] <= intermediate[4095+3569:0+3569] + a; end
12'd3570: begin if(a[3570]==1) 
	 		intermediate[4095+3570:0+3570] <= intermediate[4095+3570:0+3570] + a; end
12'd3571: begin if(a[3571]==1) 
	 		intermediate[4095+3571:0+3571] <= intermediate[4095+3571:0+3571] + a; end
12'd3572: begin if(a[3572]==1) 
	 		intermediate[4095+3572:0+3572] <= intermediate[4095+3572:0+3572] + a; end
12'd3573: begin if(a[3573]==1) 
	 		intermediate[4095+3573:0+3573] <= intermediate[4095+3573:0+3573] + a; end
12'd3574: begin if(a[3574]==1) 
	 		intermediate[4095+3574:0+3574] <= intermediate[4095+3574:0+3574] + a; end
12'd3575: begin if(a[3575]==1) 
	 		intermediate[4095+3575:0+3575] <= intermediate[4095+3575:0+3575] + a; end
12'd3576: begin if(a[3576]==1) 
	 		intermediate[4095+3576:0+3576] <= intermediate[4095+3576:0+3576] + a; end
12'd3577: begin if(a[3577]==1) 
	 		intermediate[4095+3577:0+3577] <= intermediate[4095+3577:0+3577] + a; end
12'd3578: begin if(a[3578]==1) 
	 		intermediate[4095+3578:0+3578] <= intermediate[4095+3578:0+3578] + a; end
12'd3579: begin if(a[3579]==1) 
	 		intermediate[4095+3579:0+3579] <= intermediate[4095+3579:0+3579] + a; end
12'd3580: begin if(a[3580]==1) 
	 		intermediate[4095+3580:0+3580] <= intermediate[4095+3580:0+3580] + a; end
12'd3581: begin if(a[3581]==1) 
	 		intermediate[4095+3581:0+3581] <= intermediate[4095+3581:0+3581] + a; end
12'd3582: begin if(a[3582]==1) 
	 		intermediate[4095+3582:0+3582] <= intermediate[4095+3582:0+3582] + a; end
12'd3583: begin if(a[3583]==1) 
	 		intermediate[4095+3583:0+3583] <= intermediate[4095+3583:0+3583] + a; end
12'd3584: begin if(a[3584]==1) 
	 		intermediate[4095+3584:0+3584] <= intermediate[4095+3584:0+3584] + a; end
12'd3585: begin if(a[3585]==1) 
	 		intermediate[4095+3585:0+3585] <= intermediate[4095+3585:0+3585] + a; end
12'd3586: begin if(a[3586]==1) 
	 		intermediate[4095+3586:0+3586] <= intermediate[4095+3586:0+3586] + a; end
12'd3587: begin if(a[3587]==1) 
	 		intermediate[4095+3587:0+3587] <= intermediate[4095+3587:0+3587] + a; end
12'd3588: begin if(a[3588]==1) 
	 		intermediate[4095+3588:0+3588] <= intermediate[4095+3588:0+3588] + a; end
12'd3589: begin if(a[3589]==1) 
	 		intermediate[4095+3589:0+3589] <= intermediate[4095+3589:0+3589] + a; end
12'd3590: begin if(a[3590]==1) 
	 		intermediate[4095+3590:0+3590] <= intermediate[4095+3590:0+3590] + a; end
12'd3591: begin if(a[3591]==1) 
	 		intermediate[4095+3591:0+3591] <= intermediate[4095+3591:0+3591] + a; end
12'd3592: begin if(a[3592]==1) 
	 		intermediate[4095+3592:0+3592] <= intermediate[4095+3592:0+3592] + a; end
12'd3593: begin if(a[3593]==1) 
	 		intermediate[4095+3593:0+3593] <= intermediate[4095+3593:0+3593] + a; end
12'd3594: begin if(a[3594]==1) 
	 		intermediate[4095+3594:0+3594] <= intermediate[4095+3594:0+3594] + a; end
12'd3595: begin if(a[3595]==1) 
	 		intermediate[4095+3595:0+3595] <= intermediate[4095+3595:0+3595] + a; end
12'd3596: begin if(a[3596]==1) 
	 		intermediate[4095+3596:0+3596] <= intermediate[4095+3596:0+3596] + a; end
12'd3597: begin if(a[3597]==1) 
	 		intermediate[4095+3597:0+3597] <= intermediate[4095+3597:0+3597] + a; end
12'd3598: begin if(a[3598]==1) 
	 		intermediate[4095+3598:0+3598] <= intermediate[4095+3598:0+3598] + a; end
12'd3599: begin if(a[3599]==1) 
	 		intermediate[4095+3599:0+3599] <= intermediate[4095+3599:0+3599] + a; end
12'd3600: begin if(a[3600]==1) 
	 		intermediate[4095+3600:0+3600] <= intermediate[4095+3600:0+3600] + a; end
12'd3601: begin if(a[3601]==1) 
	 		intermediate[4095+3601:0+3601] <= intermediate[4095+3601:0+3601] + a; end
12'd3602: begin if(a[3602]==1) 
	 		intermediate[4095+3602:0+3602] <= intermediate[4095+3602:0+3602] + a; end
12'd3603: begin if(a[3603]==1) 
	 		intermediate[4095+3603:0+3603] <= intermediate[4095+3603:0+3603] + a; end
12'd3604: begin if(a[3604]==1) 
	 		intermediate[4095+3604:0+3604] <= intermediate[4095+3604:0+3604] + a; end
12'd3605: begin if(a[3605]==1) 
	 		intermediate[4095+3605:0+3605] <= intermediate[4095+3605:0+3605] + a; end
12'd3606: begin if(a[3606]==1) 
	 		intermediate[4095+3606:0+3606] <= intermediate[4095+3606:0+3606] + a; end
12'd3607: begin if(a[3607]==1) 
	 		intermediate[4095+3607:0+3607] <= intermediate[4095+3607:0+3607] + a; end
12'd3608: begin if(a[3608]==1) 
	 		intermediate[4095+3608:0+3608] <= intermediate[4095+3608:0+3608] + a; end
12'd3609: begin if(a[3609]==1) 
	 		intermediate[4095+3609:0+3609] <= intermediate[4095+3609:0+3609] + a; end
12'd3610: begin if(a[3610]==1) 
	 		intermediate[4095+3610:0+3610] <= intermediate[4095+3610:0+3610] + a; end
12'd3611: begin if(a[3611]==1) 
	 		intermediate[4095+3611:0+3611] <= intermediate[4095+3611:0+3611] + a; end
12'd3612: begin if(a[3612]==1) 
	 		intermediate[4095+3612:0+3612] <= intermediate[4095+3612:0+3612] + a; end
12'd3613: begin if(a[3613]==1) 
	 		intermediate[4095+3613:0+3613] <= intermediate[4095+3613:0+3613] + a; end
12'd3614: begin if(a[3614]==1) 
	 		intermediate[4095+3614:0+3614] <= intermediate[4095+3614:0+3614] + a; end
12'd3615: begin if(a[3615]==1) 
	 		intermediate[4095+3615:0+3615] <= intermediate[4095+3615:0+3615] + a; end
12'd3616: begin if(a[3616]==1) 
	 		intermediate[4095+3616:0+3616] <= intermediate[4095+3616:0+3616] + a; end
12'd3617: begin if(a[3617]==1) 
	 		intermediate[4095+3617:0+3617] <= intermediate[4095+3617:0+3617] + a; end
12'd3618: begin if(a[3618]==1) 
	 		intermediate[4095+3618:0+3618] <= intermediate[4095+3618:0+3618] + a; end
12'd3619: begin if(a[3619]==1) 
	 		intermediate[4095+3619:0+3619] <= intermediate[4095+3619:0+3619] + a; end
12'd3620: begin if(a[3620]==1) 
	 		intermediate[4095+3620:0+3620] <= intermediate[4095+3620:0+3620] + a; end
12'd3621: begin if(a[3621]==1) 
	 		intermediate[4095+3621:0+3621] <= intermediate[4095+3621:0+3621] + a; end
12'd3622: begin if(a[3622]==1) 
	 		intermediate[4095+3622:0+3622] <= intermediate[4095+3622:0+3622] + a; end
12'd3623: begin if(a[3623]==1) 
	 		intermediate[4095+3623:0+3623] <= intermediate[4095+3623:0+3623] + a; end
12'd3624: begin if(a[3624]==1) 
	 		intermediate[4095+3624:0+3624] <= intermediate[4095+3624:0+3624] + a; end
12'd3625: begin if(a[3625]==1) 
	 		intermediate[4095+3625:0+3625] <= intermediate[4095+3625:0+3625] + a; end
12'd3626: begin if(a[3626]==1) 
	 		intermediate[4095+3626:0+3626] <= intermediate[4095+3626:0+3626] + a; end
12'd3627: begin if(a[3627]==1) 
	 		intermediate[4095+3627:0+3627] <= intermediate[4095+3627:0+3627] + a; end
12'd3628: begin if(a[3628]==1) 
	 		intermediate[4095+3628:0+3628] <= intermediate[4095+3628:0+3628] + a; end
12'd3629: begin if(a[3629]==1) 
	 		intermediate[4095+3629:0+3629] <= intermediate[4095+3629:0+3629] + a; end
12'd3630: begin if(a[3630]==1) 
	 		intermediate[4095+3630:0+3630] <= intermediate[4095+3630:0+3630] + a; end
12'd3631: begin if(a[3631]==1) 
	 		intermediate[4095+3631:0+3631] <= intermediate[4095+3631:0+3631] + a; end
12'd3632: begin if(a[3632]==1) 
	 		intermediate[4095+3632:0+3632] <= intermediate[4095+3632:0+3632] + a; end
12'd3633: begin if(a[3633]==1) 
	 		intermediate[4095+3633:0+3633] <= intermediate[4095+3633:0+3633] + a; end
12'd3634: begin if(a[3634]==1) 
	 		intermediate[4095+3634:0+3634] <= intermediate[4095+3634:0+3634] + a; end
12'd3635: begin if(a[3635]==1) 
	 		intermediate[4095+3635:0+3635] <= intermediate[4095+3635:0+3635] + a; end
12'd3636: begin if(a[3636]==1) 
	 		intermediate[4095+3636:0+3636] <= intermediate[4095+3636:0+3636] + a; end
12'd3637: begin if(a[3637]==1) 
	 		intermediate[4095+3637:0+3637] <= intermediate[4095+3637:0+3637] + a; end
12'd3638: begin if(a[3638]==1) 
	 		intermediate[4095+3638:0+3638] <= intermediate[4095+3638:0+3638] + a; end
12'd3639: begin if(a[3639]==1) 
	 		intermediate[4095+3639:0+3639] <= intermediate[4095+3639:0+3639] + a; end
12'd3640: begin if(a[3640]==1) 
	 		intermediate[4095+3640:0+3640] <= intermediate[4095+3640:0+3640] + a; end
12'd3641: begin if(a[3641]==1) 
	 		intermediate[4095+3641:0+3641] <= intermediate[4095+3641:0+3641] + a; end
12'd3642: begin if(a[3642]==1) 
	 		intermediate[4095+3642:0+3642] <= intermediate[4095+3642:0+3642] + a; end
12'd3643: begin if(a[3643]==1) 
	 		intermediate[4095+3643:0+3643] <= intermediate[4095+3643:0+3643] + a; end
12'd3644: begin if(a[3644]==1) 
	 		intermediate[4095+3644:0+3644] <= intermediate[4095+3644:0+3644] + a; end
12'd3645: begin if(a[3645]==1) 
	 		intermediate[4095+3645:0+3645] <= intermediate[4095+3645:0+3645] + a; end
12'd3646: begin if(a[3646]==1) 
	 		intermediate[4095+3646:0+3646] <= intermediate[4095+3646:0+3646] + a; end
12'd3647: begin if(a[3647]==1) 
	 		intermediate[4095+3647:0+3647] <= intermediate[4095+3647:0+3647] + a; end
12'd3648: begin if(a[3648]==1) 
	 		intermediate[4095+3648:0+3648] <= intermediate[4095+3648:0+3648] + a; end
12'd3649: begin if(a[3649]==1) 
	 		intermediate[4095+3649:0+3649] <= intermediate[4095+3649:0+3649] + a; end
12'd3650: begin if(a[3650]==1) 
	 		intermediate[4095+3650:0+3650] <= intermediate[4095+3650:0+3650] + a; end
12'd3651: begin if(a[3651]==1) 
	 		intermediate[4095+3651:0+3651] <= intermediate[4095+3651:0+3651] + a; end
12'd3652: begin if(a[3652]==1) 
	 		intermediate[4095+3652:0+3652] <= intermediate[4095+3652:0+3652] + a; end
12'd3653: begin if(a[3653]==1) 
	 		intermediate[4095+3653:0+3653] <= intermediate[4095+3653:0+3653] + a; end
12'd3654: begin if(a[3654]==1) 
	 		intermediate[4095+3654:0+3654] <= intermediate[4095+3654:0+3654] + a; end
12'd3655: begin if(a[3655]==1) 
	 		intermediate[4095+3655:0+3655] <= intermediate[4095+3655:0+3655] + a; end
12'd3656: begin if(a[3656]==1) 
	 		intermediate[4095+3656:0+3656] <= intermediate[4095+3656:0+3656] + a; end
12'd3657: begin if(a[3657]==1) 
	 		intermediate[4095+3657:0+3657] <= intermediate[4095+3657:0+3657] + a; end
12'd3658: begin if(a[3658]==1) 
	 		intermediate[4095+3658:0+3658] <= intermediate[4095+3658:0+3658] + a; end
12'd3659: begin if(a[3659]==1) 
	 		intermediate[4095+3659:0+3659] <= intermediate[4095+3659:0+3659] + a; end
12'd3660: begin if(a[3660]==1) 
	 		intermediate[4095+3660:0+3660] <= intermediate[4095+3660:0+3660] + a; end
12'd3661: begin if(a[3661]==1) 
	 		intermediate[4095+3661:0+3661] <= intermediate[4095+3661:0+3661] + a; end
12'd3662: begin if(a[3662]==1) 
	 		intermediate[4095+3662:0+3662] <= intermediate[4095+3662:0+3662] + a; end
12'd3663: begin if(a[3663]==1) 
	 		intermediate[4095+3663:0+3663] <= intermediate[4095+3663:0+3663] + a; end
12'd3664: begin if(a[3664]==1) 
	 		intermediate[4095+3664:0+3664] <= intermediate[4095+3664:0+3664] + a; end
12'd3665: begin if(a[3665]==1) 
	 		intermediate[4095+3665:0+3665] <= intermediate[4095+3665:0+3665] + a; end
12'd3666: begin if(a[3666]==1) 
	 		intermediate[4095+3666:0+3666] <= intermediate[4095+3666:0+3666] + a; end
12'd3667: begin if(a[3667]==1) 
	 		intermediate[4095+3667:0+3667] <= intermediate[4095+3667:0+3667] + a; end
12'd3668: begin if(a[3668]==1) 
	 		intermediate[4095+3668:0+3668] <= intermediate[4095+3668:0+3668] + a; end
12'd3669: begin if(a[3669]==1) 
	 		intermediate[4095+3669:0+3669] <= intermediate[4095+3669:0+3669] + a; end
12'd3670: begin if(a[3670]==1) 
	 		intermediate[4095+3670:0+3670] <= intermediate[4095+3670:0+3670] + a; end
12'd3671: begin if(a[3671]==1) 
	 		intermediate[4095+3671:0+3671] <= intermediate[4095+3671:0+3671] + a; end
12'd3672: begin if(a[3672]==1) 
	 		intermediate[4095+3672:0+3672] <= intermediate[4095+3672:0+3672] + a; end
12'd3673: begin if(a[3673]==1) 
	 		intermediate[4095+3673:0+3673] <= intermediate[4095+3673:0+3673] + a; end
12'd3674: begin if(a[3674]==1) 
	 		intermediate[4095+3674:0+3674] <= intermediate[4095+3674:0+3674] + a; end
12'd3675: begin if(a[3675]==1) 
	 		intermediate[4095+3675:0+3675] <= intermediate[4095+3675:0+3675] + a; end
12'd3676: begin if(a[3676]==1) 
	 		intermediate[4095+3676:0+3676] <= intermediate[4095+3676:0+3676] + a; end
12'd3677: begin if(a[3677]==1) 
	 		intermediate[4095+3677:0+3677] <= intermediate[4095+3677:0+3677] + a; end
12'd3678: begin if(a[3678]==1) 
	 		intermediate[4095+3678:0+3678] <= intermediate[4095+3678:0+3678] + a; end
12'd3679: begin if(a[3679]==1) 
	 		intermediate[4095+3679:0+3679] <= intermediate[4095+3679:0+3679] + a; end
12'd3680: begin if(a[3680]==1) 
	 		intermediate[4095+3680:0+3680] <= intermediate[4095+3680:0+3680] + a; end
12'd3681: begin if(a[3681]==1) 
	 		intermediate[4095+3681:0+3681] <= intermediate[4095+3681:0+3681] + a; end
12'd3682: begin if(a[3682]==1) 
	 		intermediate[4095+3682:0+3682] <= intermediate[4095+3682:0+3682] + a; end
12'd3683: begin if(a[3683]==1) 
	 		intermediate[4095+3683:0+3683] <= intermediate[4095+3683:0+3683] + a; end
12'd3684: begin if(a[3684]==1) 
	 		intermediate[4095+3684:0+3684] <= intermediate[4095+3684:0+3684] + a; end
12'd3685: begin if(a[3685]==1) 
	 		intermediate[4095+3685:0+3685] <= intermediate[4095+3685:0+3685] + a; end
12'd3686: begin if(a[3686]==1) 
	 		intermediate[4095+3686:0+3686] <= intermediate[4095+3686:0+3686] + a; end
12'd3687: begin if(a[3687]==1) 
	 		intermediate[4095+3687:0+3687] <= intermediate[4095+3687:0+3687] + a; end
12'd3688: begin if(a[3688]==1) 
	 		intermediate[4095+3688:0+3688] <= intermediate[4095+3688:0+3688] + a; end
12'd3689: begin if(a[3689]==1) 
	 		intermediate[4095+3689:0+3689] <= intermediate[4095+3689:0+3689] + a; end
12'd3690: begin if(a[3690]==1) 
	 		intermediate[4095+3690:0+3690] <= intermediate[4095+3690:0+3690] + a; end
12'd3691: begin if(a[3691]==1) 
	 		intermediate[4095+3691:0+3691] <= intermediate[4095+3691:0+3691] + a; end
12'd3692: begin if(a[3692]==1) 
	 		intermediate[4095+3692:0+3692] <= intermediate[4095+3692:0+3692] + a; end
12'd3693: begin if(a[3693]==1) 
	 		intermediate[4095+3693:0+3693] <= intermediate[4095+3693:0+3693] + a; end
12'd3694: begin if(a[3694]==1) 
	 		intermediate[4095+3694:0+3694] <= intermediate[4095+3694:0+3694] + a; end
12'd3695: begin if(a[3695]==1) 
	 		intermediate[4095+3695:0+3695] <= intermediate[4095+3695:0+3695] + a; end
12'd3696: begin if(a[3696]==1) 
	 		intermediate[4095+3696:0+3696] <= intermediate[4095+3696:0+3696] + a; end
12'd3697: begin if(a[3697]==1) 
	 		intermediate[4095+3697:0+3697] <= intermediate[4095+3697:0+3697] + a; end
12'd3698: begin if(a[3698]==1) 
	 		intermediate[4095+3698:0+3698] <= intermediate[4095+3698:0+3698] + a; end
12'd3699: begin if(a[3699]==1) 
	 		intermediate[4095+3699:0+3699] <= intermediate[4095+3699:0+3699] + a; end
12'd3700: begin if(a[3700]==1) 
	 		intermediate[4095+3700:0+3700] <= intermediate[4095+3700:0+3700] + a; end
12'd3701: begin if(a[3701]==1) 
	 		intermediate[4095+3701:0+3701] <= intermediate[4095+3701:0+3701] + a; end
12'd3702: begin if(a[3702]==1) 
	 		intermediate[4095+3702:0+3702] <= intermediate[4095+3702:0+3702] + a; end
12'd3703: begin if(a[3703]==1) 
	 		intermediate[4095+3703:0+3703] <= intermediate[4095+3703:0+3703] + a; end
12'd3704: begin if(a[3704]==1) 
	 		intermediate[4095+3704:0+3704] <= intermediate[4095+3704:0+3704] + a; end
12'd3705: begin if(a[3705]==1) 
	 		intermediate[4095+3705:0+3705] <= intermediate[4095+3705:0+3705] + a; end
12'd3706: begin if(a[3706]==1) 
	 		intermediate[4095+3706:0+3706] <= intermediate[4095+3706:0+3706] + a; end
12'd3707: begin if(a[3707]==1) 
	 		intermediate[4095+3707:0+3707] <= intermediate[4095+3707:0+3707] + a; end
12'd3708: begin if(a[3708]==1) 
	 		intermediate[4095+3708:0+3708] <= intermediate[4095+3708:0+3708] + a; end
12'd3709: begin if(a[3709]==1) 
	 		intermediate[4095+3709:0+3709] <= intermediate[4095+3709:0+3709] + a; end
12'd3710: begin if(a[3710]==1) 
	 		intermediate[4095+3710:0+3710] <= intermediate[4095+3710:0+3710] + a; end
12'd3711: begin if(a[3711]==1) 
	 		intermediate[4095+3711:0+3711] <= intermediate[4095+3711:0+3711] + a; end
12'd3712: begin if(a[3712]==1) 
	 		intermediate[4095+3712:0+3712] <= intermediate[4095+3712:0+3712] + a; end
12'd3713: begin if(a[3713]==1) 
	 		intermediate[4095+3713:0+3713] <= intermediate[4095+3713:0+3713] + a; end
12'd3714: begin if(a[3714]==1) 
	 		intermediate[4095+3714:0+3714] <= intermediate[4095+3714:0+3714] + a; end
12'd3715: begin if(a[3715]==1) 
	 		intermediate[4095+3715:0+3715] <= intermediate[4095+3715:0+3715] + a; end
12'd3716: begin if(a[3716]==1) 
	 		intermediate[4095+3716:0+3716] <= intermediate[4095+3716:0+3716] + a; end
12'd3717: begin if(a[3717]==1) 
	 		intermediate[4095+3717:0+3717] <= intermediate[4095+3717:0+3717] + a; end
12'd3718: begin if(a[3718]==1) 
	 		intermediate[4095+3718:0+3718] <= intermediate[4095+3718:0+3718] + a; end
12'd3719: begin if(a[3719]==1) 
	 		intermediate[4095+3719:0+3719] <= intermediate[4095+3719:0+3719] + a; end
12'd3720: begin if(a[3720]==1) 
	 		intermediate[4095+3720:0+3720] <= intermediate[4095+3720:0+3720] + a; end
12'd3721: begin if(a[3721]==1) 
	 		intermediate[4095+3721:0+3721] <= intermediate[4095+3721:0+3721] + a; end
12'd3722: begin if(a[3722]==1) 
	 		intermediate[4095+3722:0+3722] <= intermediate[4095+3722:0+3722] + a; end
12'd3723: begin if(a[3723]==1) 
	 		intermediate[4095+3723:0+3723] <= intermediate[4095+3723:0+3723] + a; end
12'd3724: begin if(a[3724]==1) 
	 		intermediate[4095+3724:0+3724] <= intermediate[4095+3724:0+3724] + a; end
12'd3725: begin if(a[3725]==1) 
	 		intermediate[4095+3725:0+3725] <= intermediate[4095+3725:0+3725] + a; end
12'd3726: begin if(a[3726]==1) 
	 		intermediate[4095+3726:0+3726] <= intermediate[4095+3726:0+3726] + a; end
12'd3727: begin if(a[3727]==1) 
	 		intermediate[4095+3727:0+3727] <= intermediate[4095+3727:0+3727] + a; end
12'd3728: begin if(a[3728]==1) 
	 		intermediate[4095+3728:0+3728] <= intermediate[4095+3728:0+3728] + a; end
12'd3729: begin if(a[3729]==1) 
	 		intermediate[4095+3729:0+3729] <= intermediate[4095+3729:0+3729] + a; end
12'd3730: begin if(a[3730]==1) 
	 		intermediate[4095+3730:0+3730] <= intermediate[4095+3730:0+3730] + a; end
12'd3731: begin if(a[3731]==1) 
	 		intermediate[4095+3731:0+3731] <= intermediate[4095+3731:0+3731] + a; end
12'd3732: begin if(a[3732]==1) 
	 		intermediate[4095+3732:0+3732] <= intermediate[4095+3732:0+3732] + a; end
12'd3733: begin if(a[3733]==1) 
	 		intermediate[4095+3733:0+3733] <= intermediate[4095+3733:0+3733] + a; end
12'd3734: begin if(a[3734]==1) 
	 		intermediate[4095+3734:0+3734] <= intermediate[4095+3734:0+3734] + a; end
12'd3735: begin if(a[3735]==1) 
	 		intermediate[4095+3735:0+3735] <= intermediate[4095+3735:0+3735] + a; end
12'd3736: begin if(a[3736]==1) 
	 		intermediate[4095+3736:0+3736] <= intermediate[4095+3736:0+3736] + a; end
12'd3737: begin if(a[3737]==1) 
	 		intermediate[4095+3737:0+3737] <= intermediate[4095+3737:0+3737] + a; end
12'd3738: begin if(a[3738]==1) 
	 		intermediate[4095+3738:0+3738] <= intermediate[4095+3738:0+3738] + a; end
12'd3739: begin if(a[3739]==1) 
	 		intermediate[4095+3739:0+3739] <= intermediate[4095+3739:0+3739] + a; end
12'd3740: begin if(a[3740]==1) 
	 		intermediate[4095+3740:0+3740] <= intermediate[4095+3740:0+3740] + a; end
12'd3741: begin if(a[3741]==1) 
	 		intermediate[4095+3741:0+3741] <= intermediate[4095+3741:0+3741] + a; end
12'd3742: begin if(a[3742]==1) 
	 		intermediate[4095+3742:0+3742] <= intermediate[4095+3742:0+3742] + a; end
12'd3743: begin if(a[3743]==1) 
	 		intermediate[4095+3743:0+3743] <= intermediate[4095+3743:0+3743] + a; end
12'd3744: begin if(a[3744]==1) 
	 		intermediate[4095+3744:0+3744] <= intermediate[4095+3744:0+3744] + a; end
12'd3745: begin if(a[3745]==1) 
	 		intermediate[4095+3745:0+3745] <= intermediate[4095+3745:0+3745] + a; end
12'd3746: begin if(a[3746]==1) 
	 		intermediate[4095+3746:0+3746] <= intermediate[4095+3746:0+3746] + a; end
12'd3747: begin if(a[3747]==1) 
	 		intermediate[4095+3747:0+3747] <= intermediate[4095+3747:0+3747] + a; end
12'd3748: begin if(a[3748]==1) 
	 		intermediate[4095+3748:0+3748] <= intermediate[4095+3748:0+3748] + a; end
12'd3749: begin if(a[3749]==1) 
	 		intermediate[4095+3749:0+3749] <= intermediate[4095+3749:0+3749] + a; end
12'd3750: begin if(a[3750]==1) 
	 		intermediate[4095+3750:0+3750] <= intermediate[4095+3750:0+3750] + a; end
12'd3751: begin if(a[3751]==1) 
	 		intermediate[4095+3751:0+3751] <= intermediate[4095+3751:0+3751] + a; end
12'd3752: begin if(a[3752]==1) 
	 		intermediate[4095+3752:0+3752] <= intermediate[4095+3752:0+3752] + a; end
12'd3753: begin if(a[3753]==1) 
	 		intermediate[4095+3753:0+3753] <= intermediate[4095+3753:0+3753] + a; end
12'd3754: begin if(a[3754]==1) 
	 		intermediate[4095+3754:0+3754] <= intermediate[4095+3754:0+3754] + a; end
12'd3755: begin if(a[3755]==1) 
	 		intermediate[4095+3755:0+3755] <= intermediate[4095+3755:0+3755] + a; end
12'd3756: begin if(a[3756]==1) 
	 		intermediate[4095+3756:0+3756] <= intermediate[4095+3756:0+3756] + a; end
12'd3757: begin if(a[3757]==1) 
	 		intermediate[4095+3757:0+3757] <= intermediate[4095+3757:0+3757] + a; end
12'd3758: begin if(a[3758]==1) 
	 		intermediate[4095+3758:0+3758] <= intermediate[4095+3758:0+3758] + a; end
12'd3759: begin if(a[3759]==1) 
	 		intermediate[4095+3759:0+3759] <= intermediate[4095+3759:0+3759] + a; end
12'd3760: begin if(a[3760]==1) 
	 		intermediate[4095+3760:0+3760] <= intermediate[4095+3760:0+3760] + a; end
12'd3761: begin if(a[3761]==1) 
	 		intermediate[4095+3761:0+3761] <= intermediate[4095+3761:0+3761] + a; end
12'd3762: begin if(a[3762]==1) 
	 		intermediate[4095+3762:0+3762] <= intermediate[4095+3762:0+3762] + a; end
12'd3763: begin if(a[3763]==1) 
	 		intermediate[4095+3763:0+3763] <= intermediate[4095+3763:0+3763] + a; end
12'd3764: begin if(a[3764]==1) 
	 		intermediate[4095+3764:0+3764] <= intermediate[4095+3764:0+3764] + a; end
12'd3765: begin if(a[3765]==1) 
	 		intermediate[4095+3765:0+3765] <= intermediate[4095+3765:0+3765] + a; end
12'd3766: begin if(a[3766]==1) 
	 		intermediate[4095+3766:0+3766] <= intermediate[4095+3766:0+3766] + a; end
12'd3767: begin if(a[3767]==1) 
	 		intermediate[4095+3767:0+3767] <= intermediate[4095+3767:0+3767] + a; end
12'd3768: begin if(a[3768]==1) 
	 		intermediate[4095+3768:0+3768] <= intermediate[4095+3768:0+3768] + a; end
12'd3769: begin if(a[3769]==1) 
	 		intermediate[4095+3769:0+3769] <= intermediate[4095+3769:0+3769] + a; end
12'd3770: begin if(a[3770]==1) 
	 		intermediate[4095+3770:0+3770] <= intermediate[4095+3770:0+3770] + a; end
12'd3771: begin if(a[3771]==1) 
	 		intermediate[4095+3771:0+3771] <= intermediate[4095+3771:0+3771] + a; end
12'd3772: begin if(a[3772]==1) 
	 		intermediate[4095+3772:0+3772] <= intermediate[4095+3772:0+3772] + a; end
12'd3773: begin if(a[3773]==1) 
	 		intermediate[4095+3773:0+3773] <= intermediate[4095+3773:0+3773] + a; end
12'd3774: begin if(a[3774]==1) 
	 		intermediate[4095+3774:0+3774] <= intermediate[4095+3774:0+3774] + a; end
12'd3775: begin if(a[3775]==1) 
	 		intermediate[4095+3775:0+3775] <= intermediate[4095+3775:0+3775] + a; end
12'd3776: begin if(a[3776]==1) 
	 		intermediate[4095+3776:0+3776] <= intermediate[4095+3776:0+3776] + a; end
12'd3777: begin if(a[3777]==1) 
	 		intermediate[4095+3777:0+3777] <= intermediate[4095+3777:0+3777] + a; end
12'd3778: begin if(a[3778]==1) 
	 		intermediate[4095+3778:0+3778] <= intermediate[4095+3778:0+3778] + a; end
12'd3779: begin if(a[3779]==1) 
	 		intermediate[4095+3779:0+3779] <= intermediate[4095+3779:0+3779] + a; end
12'd3780: begin if(a[3780]==1) 
	 		intermediate[4095+3780:0+3780] <= intermediate[4095+3780:0+3780] + a; end
12'd3781: begin if(a[3781]==1) 
	 		intermediate[4095+3781:0+3781] <= intermediate[4095+3781:0+3781] + a; end
12'd3782: begin if(a[3782]==1) 
	 		intermediate[4095+3782:0+3782] <= intermediate[4095+3782:0+3782] + a; end
12'd3783: begin if(a[3783]==1) 
	 		intermediate[4095+3783:0+3783] <= intermediate[4095+3783:0+3783] + a; end
12'd3784: begin if(a[3784]==1) 
	 		intermediate[4095+3784:0+3784] <= intermediate[4095+3784:0+3784] + a; end
12'd3785: begin if(a[3785]==1) 
	 		intermediate[4095+3785:0+3785] <= intermediate[4095+3785:0+3785] + a; end
12'd3786: begin if(a[3786]==1) 
	 		intermediate[4095+3786:0+3786] <= intermediate[4095+3786:0+3786] + a; end
12'd3787: begin if(a[3787]==1) 
	 		intermediate[4095+3787:0+3787] <= intermediate[4095+3787:0+3787] + a; end
12'd3788: begin if(a[3788]==1) 
	 		intermediate[4095+3788:0+3788] <= intermediate[4095+3788:0+3788] + a; end
12'd3789: begin if(a[3789]==1) 
	 		intermediate[4095+3789:0+3789] <= intermediate[4095+3789:0+3789] + a; end
12'd3790: begin if(a[3790]==1) 
	 		intermediate[4095+3790:0+3790] <= intermediate[4095+3790:0+3790] + a; end
12'd3791: begin if(a[3791]==1) 
	 		intermediate[4095+3791:0+3791] <= intermediate[4095+3791:0+3791] + a; end
12'd3792: begin if(a[3792]==1) 
	 		intermediate[4095+3792:0+3792] <= intermediate[4095+3792:0+3792] + a; end
12'd3793: begin if(a[3793]==1) 
	 		intermediate[4095+3793:0+3793] <= intermediate[4095+3793:0+3793] + a; end
12'd3794: begin if(a[3794]==1) 
	 		intermediate[4095+3794:0+3794] <= intermediate[4095+3794:0+3794] + a; end
12'd3795: begin if(a[3795]==1) 
	 		intermediate[4095+3795:0+3795] <= intermediate[4095+3795:0+3795] + a; end
12'd3796: begin if(a[3796]==1) 
	 		intermediate[4095+3796:0+3796] <= intermediate[4095+3796:0+3796] + a; end
12'd3797: begin if(a[3797]==1) 
	 		intermediate[4095+3797:0+3797] <= intermediate[4095+3797:0+3797] + a; end
12'd3798: begin if(a[3798]==1) 
	 		intermediate[4095+3798:0+3798] <= intermediate[4095+3798:0+3798] + a; end
12'd3799: begin if(a[3799]==1) 
	 		intermediate[4095+3799:0+3799] <= intermediate[4095+3799:0+3799] + a; end
12'd3800: begin if(a[3800]==1) 
	 		intermediate[4095+3800:0+3800] <= intermediate[4095+3800:0+3800] + a; end
12'd3801: begin if(a[3801]==1) 
	 		intermediate[4095+3801:0+3801] <= intermediate[4095+3801:0+3801] + a; end
12'd3802: begin if(a[3802]==1) 
	 		intermediate[4095+3802:0+3802] <= intermediate[4095+3802:0+3802] + a; end
12'd3803: begin if(a[3803]==1) 
	 		intermediate[4095+3803:0+3803] <= intermediate[4095+3803:0+3803] + a; end
12'd3804: begin if(a[3804]==1) 
	 		intermediate[4095+3804:0+3804] <= intermediate[4095+3804:0+3804] + a; end
12'd3805: begin if(a[3805]==1) 
	 		intermediate[4095+3805:0+3805] <= intermediate[4095+3805:0+3805] + a; end
12'd3806: begin if(a[3806]==1) 
	 		intermediate[4095+3806:0+3806] <= intermediate[4095+3806:0+3806] + a; end
12'd3807: begin if(a[3807]==1) 
	 		intermediate[4095+3807:0+3807] <= intermediate[4095+3807:0+3807] + a; end
12'd3808: begin if(a[3808]==1) 
	 		intermediate[4095+3808:0+3808] <= intermediate[4095+3808:0+3808] + a; end
12'd3809: begin if(a[3809]==1) 
	 		intermediate[4095+3809:0+3809] <= intermediate[4095+3809:0+3809] + a; end
12'd3810: begin if(a[3810]==1) 
	 		intermediate[4095+3810:0+3810] <= intermediate[4095+3810:0+3810] + a; end
12'd3811: begin if(a[3811]==1) 
	 		intermediate[4095+3811:0+3811] <= intermediate[4095+3811:0+3811] + a; end
12'd3812: begin if(a[3812]==1) 
	 		intermediate[4095+3812:0+3812] <= intermediate[4095+3812:0+3812] + a; end
12'd3813: begin if(a[3813]==1) 
	 		intermediate[4095+3813:0+3813] <= intermediate[4095+3813:0+3813] + a; end
12'd3814: begin if(a[3814]==1) 
	 		intermediate[4095+3814:0+3814] <= intermediate[4095+3814:0+3814] + a; end
12'd3815: begin if(a[3815]==1) 
	 		intermediate[4095+3815:0+3815] <= intermediate[4095+3815:0+3815] + a; end
12'd3816: begin if(a[3816]==1) 
	 		intermediate[4095+3816:0+3816] <= intermediate[4095+3816:0+3816] + a; end
12'd3817: begin if(a[3817]==1) 
	 		intermediate[4095+3817:0+3817] <= intermediate[4095+3817:0+3817] + a; end
12'd3818: begin if(a[3818]==1) 
	 		intermediate[4095+3818:0+3818] <= intermediate[4095+3818:0+3818] + a; end
12'd3819: begin if(a[3819]==1) 
	 		intermediate[4095+3819:0+3819] <= intermediate[4095+3819:0+3819] + a; end
12'd3820: begin if(a[3820]==1) 
	 		intermediate[4095+3820:0+3820] <= intermediate[4095+3820:0+3820] + a; end
12'd3821: begin if(a[3821]==1) 
	 		intermediate[4095+3821:0+3821] <= intermediate[4095+3821:0+3821] + a; end
12'd3822: begin if(a[3822]==1) 
	 		intermediate[4095+3822:0+3822] <= intermediate[4095+3822:0+3822] + a; end
12'd3823: begin if(a[3823]==1) 
	 		intermediate[4095+3823:0+3823] <= intermediate[4095+3823:0+3823] + a; end
12'd3824: begin if(a[3824]==1) 
	 		intermediate[4095+3824:0+3824] <= intermediate[4095+3824:0+3824] + a; end
12'd3825: begin if(a[3825]==1) 
	 		intermediate[4095+3825:0+3825] <= intermediate[4095+3825:0+3825] + a; end
12'd3826: begin if(a[3826]==1) 
	 		intermediate[4095+3826:0+3826] <= intermediate[4095+3826:0+3826] + a; end
12'd3827: begin if(a[3827]==1) 
	 		intermediate[4095+3827:0+3827] <= intermediate[4095+3827:0+3827] + a; end
12'd3828: begin if(a[3828]==1) 
	 		intermediate[4095+3828:0+3828] <= intermediate[4095+3828:0+3828] + a; end
12'd3829: begin if(a[3829]==1) 
	 		intermediate[4095+3829:0+3829] <= intermediate[4095+3829:0+3829] + a; end
12'd3830: begin if(a[3830]==1) 
	 		intermediate[4095+3830:0+3830] <= intermediate[4095+3830:0+3830] + a; end
12'd3831: begin if(a[3831]==1) 
	 		intermediate[4095+3831:0+3831] <= intermediate[4095+3831:0+3831] + a; end
12'd3832: begin if(a[3832]==1) 
	 		intermediate[4095+3832:0+3832] <= intermediate[4095+3832:0+3832] + a; end
12'd3833: begin if(a[3833]==1) 
	 		intermediate[4095+3833:0+3833] <= intermediate[4095+3833:0+3833] + a; end
12'd3834: begin if(a[3834]==1) 
	 		intermediate[4095+3834:0+3834] <= intermediate[4095+3834:0+3834] + a; end
12'd3835: begin if(a[3835]==1) 
	 		intermediate[4095+3835:0+3835] <= intermediate[4095+3835:0+3835] + a; end
12'd3836: begin if(a[3836]==1) 
	 		intermediate[4095+3836:0+3836] <= intermediate[4095+3836:0+3836] + a; end
12'd3837: begin if(a[3837]==1) 
	 		intermediate[4095+3837:0+3837] <= intermediate[4095+3837:0+3837] + a; end
12'd3838: begin if(a[3838]==1) 
	 		intermediate[4095+3838:0+3838] <= intermediate[4095+3838:0+3838] + a; end
12'd3839: begin if(a[3839]==1) 
	 		intermediate[4095+3839:0+3839] <= intermediate[4095+3839:0+3839] + a; end
12'd3840: begin if(a[3840]==1) 
	 		intermediate[4095+3840:0+3840] <= intermediate[4095+3840:0+3840] + a; end
12'd3841: begin if(a[3841]==1) 
	 		intermediate[4095+3841:0+3841] <= intermediate[4095+3841:0+3841] + a; end
12'd3842: begin if(a[3842]==1) 
	 		intermediate[4095+3842:0+3842] <= intermediate[4095+3842:0+3842] + a; end
12'd3843: begin if(a[3843]==1) 
	 		intermediate[4095+3843:0+3843] <= intermediate[4095+3843:0+3843] + a; end
12'd3844: begin if(a[3844]==1) 
	 		intermediate[4095+3844:0+3844] <= intermediate[4095+3844:0+3844] + a; end
12'd3845: begin if(a[3845]==1) 
	 		intermediate[4095+3845:0+3845] <= intermediate[4095+3845:0+3845] + a; end
12'd3846: begin if(a[3846]==1) 
	 		intermediate[4095+3846:0+3846] <= intermediate[4095+3846:0+3846] + a; end
12'd3847: begin if(a[3847]==1) 
	 		intermediate[4095+3847:0+3847] <= intermediate[4095+3847:0+3847] + a; end
12'd3848: begin if(a[3848]==1) 
	 		intermediate[4095+3848:0+3848] <= intermediate[4095+3848:0+3848] + a; end
12'd3849: begin if(a[3849]==1) 
	 		intermediate[4095+3849:0+3849] <= intermediate[4095+3849:0+3849] + a; end
12'd3850: begin if(a[3850]==1) 
	 		intermediate[4095+3850:0+3850] <= intermediate[4095+3850:0+3850] + a; end
12'd3851: begin if(a[3851]==1) 
	 		intermediate[4095+3851:0+3851] <= intermediate[4095+3851:0+3851] + a; end
12'd3852: begin if(a[3852]==1) 
	 		intermediate[4095+3852:0+3852] <= intermediate[4095+3852:0+3852] + a; end
12'd3853: begin if(a[3853]==1) 
	 		intermediate[4095+3853:0+3853] <= intermediate[4095+3853:0+3853] + a; end
12'd3854: begin if(a[3854]==1) 
	 		intermediate[4095+3854:0+3854] <= intermediate[4095+3854:0+3854] + a; end
12'd3855: begin if(a[3855]==1) 
	 		intermediate[4095+3855:0+3855] <= intermediate[4095+3855:0+3855] + a; end
12'd3856: begin if(a[3856]==1) 
	 		intermediate[4095+3856:0+3856] <= intermediate[4095+3856:0+3856] + a; end
12'd3857: begin if(a[3857]==1) 
	 		intermediate[4095+3857:0+3857] <= intermediate[4095+3857:0+3857] + a; end
12'd3858: begin if(a[3858]==1) 
	 		intermediate[4095+3858:0+3858] <= intermediate[4095+3858:0+3858] + a; end
12'd3859: begin if(a[3859]==1) 
	 		intermediate[4095+3859:0+3859] <= intermediate[4095+3859:0+3859] + a; end
12'd3860: begin if(a[3860]==1) 
	 		intermediate[4095+3860:0+3860] <= intermediate[4095+3860:0+3860] + a; end
12'd3861: begin if(a[3861]==1) 
	 		intermediate[4095+3861:0+3861] <= intermediate[4095+3861:0+3861] + a; end
12'd3862: begin if(a[3862]==1) 
	 		intermediate[4095+3862:0+3862] <= intermediate[4095+3862:0+3862] + a; end
12'd3863: begin if(a[3863]==1) 
	 		intermediate[4095+3863:0+3863] <= intermediate[4095+3863:0+3863] + a; end
12'd3864: begin if(a[3864]==1) 
	 		intermediate[4095+3864:0+3864] <= intermediate[4095+3864:0+3864] + a; end
12'd3865: begin if(a[3865]==1) 
	 		intermediate[4095+3865:0+3865] <= intermediate[4095+3865:0+3865] + a; end
12'd3866: begin if(a[3866]==1) 
	 		intermediate[4095+3866:0+3866] <= intermediate[4095+3866:0+3866] + a; end
12'd3867: begin if(a[3867]==1) 
	 		intermediate[4095+3867:0+3867] <= intermediate[4095+3867:0+3867] + a; end
12'd3868: begin if(a[3868]==1) 
	 		intermediate[4095+3868:0+3868] <= intermediate[4095+3868:0+3868] + a; end
12'd3869: begin if(a[3869]==1) 
	 		intermediate[4095+3869:0+3869] <= intermediate[4095+3869:0+3869] + a; end
12'd3870: begin if(a[3870]==1) 
	 		intermediate[4095+3870:0+3870] <= intermediate[4095+3870:0+3870] + a; end
12'd3871: begin if(a[3871]==1) 
	 		intermediate[4095+3871:0+3871] <= intermediate[4095+3871:0+3871] + a; end
12'd3872: begin if(a[3872]==1) 
	 		intermediate[4095+3872:0+3872] <= intermediate[4095+3872:0+3872] + a; end
12'd3873: begin if(a[3873]==1) 
	 		intermediate[4095+3873:0+3873] <= intermediate[4095+3873:0+3873] + a; end
12'd3874: begin if(a[3874]==1) 
	 		intermediate[4095+3874:0+3874] <= intermediate[4095+3874:0+3874] + a; end
12'd3875: begin if(a[3875]==1) 
	 		intermediate[4095+3875:0+3875] <= intermediate[4095+3875:0+3875] + a; end
12'd3876: begin if(a[3876]==1) 
	 		intermediate[4095+3876:0+3876] <= intermediate[4095+3876:0+3876] + a; end
12'd3877: begin if(a[3877]==1) 
	 		intermediate[4095+3877:0+3877] <= intermediate[4095+3877:0+3877] + a; end
12'd3878: begin if(a[3878]==1) 
	 		intermediate[4095+3878:0+3878] <= intermediate[4095+3878:0+3878] + a; end
12'd3879: begin if(a[3879]==1) 
	 		intermediate[4095+3879:0+3879] <= intermediate[4095+3879:0+3879] + a; end
12'd3880: begin if(a[3880]==1) 
	 		intermediate[4095+3880:0+3880] <= intermediate[4095+3880:0+3880] + a; end
12'd3881: begin if(a[3881]==1) 
	 		intermediate[4095+3881:0+3881] <= intermediate[4095+3881:0+3881] + a; end
12'd3882: begin if(a[3882]==1) 
	 		intermediate[4095+3882:0+3882] <= intermediate[4095+3882:0+3882] + a; end
12'd3883: begin if(a[3883]==1) 
	 		intermediate[4095+3883:0+3883] <= intermediate[4095+3883:0+3883] + a; end
12'd3884: begin if(a[3884]==1) 
	 		intermediate[4095+3884:0+3884] <= intermediate[4095+3884:0+3884] + a; end
12'd3885: begin if(a[3885]==1) 
	 		intermediate[4095+3885:0+3885] <= intermediate[4095+3885:0+3885] + a; end
12'd3886: begin if(a[3886]==1) 
	 		intermediate[4095+3886:0+3886] <= intermediate[4095+3886:0+3886] + a; end
12'd3887: begin if(a[3887]==1) 
	 		intermediate[4095+3887:0+3887] <= intermediate[4095+3887:0+3887] + a; end
12'd3888: begin if(a[3888]==1) 
	 		intermediate[4095+3888:0+3888] <= intermediate[4095+3888:0+3888] + a; end
12'd3889: begin if(a[3889]==1) 
	 		intermediate[4095+3889:0+3889] <= intermediate[4095+3889:0+3889] + a; end
12'd3890: begin if(a[3890]==1) 
	 		intermediate[4095+3890:0+3890] <= intermediate[4095+3890:0+3890] + a; end
12'd3891: begin if(a[3891]==1) 
	 		intermediate[4095+3891:0+3891] <= intermediate[4095+3891:0+3891] + a; end
12'd3892: begin if(a[3892]==1) 
	 		intermediate[4095+3892:0+3892] <= intermediate[4095+3892:0+3892] + a; end
12'd3893: begin if(a[3893]==1) 
	 		intermediate[4095+3893:0+3893] <= intermediate[4095+3893:0+3893] + a; end
12'd3894: begin if(a[3894]==1) 
	 		intermediate[4095+3894:0+3894] <= intermediate[4095+3894:0+3894] + a; end
12'd3895: begin if(a[3895]==1) 
	 		intermediate[4095+3895:0+3895] <= intermediate[4095+3895:0+3895] + a; end
12'd3896: begin if(a[3896]==1) 
	 		intermediate[4095+3896:0+3896] <= intermediate[4095+3896:0+3896] + a; end
12'd3897: begin if(a[3897]==1) 
	 		intermediate[4095+3897:0+3897] <= intermediate[4095+3897:0+3897] + a; end
12'd3898: begin if(a[3898]==1) 
	 		intermediate[4095+3898:0+3898] <= intermediate[4095+3898:0+3898] + a; end
12'd3899: begin if(a[3899]==1) 
	 		intermediate[4095+3899:0+3899] <= intermediate[4095+3899:0+3899] + a; end
12'd3900: begin if(a[3900]==1) 
	 		intermediate[4095+3900:0+3900] <= intermediate[4095+3900:0+3900] + a; end
12'd3901: begin if(a[3901]==1) 
	 		intermediate[4095+3901:0+3901] <= intermediate[4095+3901:0+3901] + a; end
12'd3902: begin if(a[3902]==1) 
	 		intermediate[4095+3902:0+3902] <= intermediate[4095+3902:0+3902] + a; end
12'd3903: begin if(a[3903]==1) 
	 		intermediate[4095+3903:0+3903] <= intermediate[4095+3903:0+3903] + a; end
12'd3904: begin if(a[3904]==1) 
	 		intermediate[4095+3904:0+3904] <= intermediate[4095+3904:0+3904] + a; end
12'd3905: begin if(a[3905]==1) 
	 		intermediate[4095+3905:0+3905] <= intermediate[4095+3905:0+3905] + a; end
12'd3906: begin if(a[3906]==1) 
	 		intermediate[4095+3906:0+3906] <= intermediate[4095+3906:0+3906] + a; end
12'd3907: begin if(a[3907]==1) 
	 		intermediate[4095+3907:0+3907] <= intermediate[4095+3907:0+3907] + a; end
12'd3908: begin if(a[3908]==1) 
	 		intermediate[4095+3908:0+3908] <= intermediate[4095+3908:0+3908] + a; end
12'd3909: begin if(a[3909]==1) 
	 		intermediate[4095+3909:0+3909] <= intermediate[4095+3909:0+3909] + a; end
12'd3910: begin if(a[3910]==1) 
	 		intermediate[4095+3910:0+3910] <= intermediate[4095+3910:0+3910] + a; end
12'd3911: begin if(a[3911]==1) 
	 		intermediate[4095+3911:0+3911] <= intermediate[4095+3911:0+3911] + a; end
12'd3912: begin if(a[3912]==1) 
	 		intermediate[4095+3912:0+3912] <= intermediate[4095+3912:0+3912] + a; end
12'd3913: begin if(a[3913]==1) 
	 		intermediate[4095+3913:0+3913] <= intermediate[4095+3913:0+3913] + a; end
12'd3914: begin if(a[3914]==1) 
	 		intermediate[4095+3914:0+3914] <= intermediate[4095+3914:0+3914] + a; end
12'd3915: begin if(a[3915]==1) 
	 		intermediate[4095+3915:0+3915] <= intermediate[4095+3915:0+3915] + a; end
12'd3916: begin if(a[3916]==1) 
	 		intermediate[4095+3916:0+3916] <= intermediate[4095+3916:0+3916] + a; end
12'd3917: begin if(a[3917]==1) 
	 		intermediate[4095+3917:0+3917] <= intermediate[4095+3917:0+3917] + a; end
12'd3918: begin if(a[3918]==1) 
	 		intermediate[4095+3918:0+3918] <= intermediate[4095+3918:0+3918] + a; end
12'd3919: begin if(a[3919]==1) 
	 		intermediate[4095+3919:0+3919] <= intermediate[4095+3919:0+3919] + a; end
12'd3920: begin if(a[3920]==1) 
	 		intermediate[4095+3920:0+3920] <= intermediate[4095+3920:0+3920] + a; end
12'd3921: begin if(a[3921]==1) 
	 		intermediate[4095+3921:0+3921] <= intermediate[4095+3921:0+3921] + a; end
12'd3922: begin if(a[3922]==1) 
	 		intermediate[4095+3922:0+3922] <= intermediate[4095+3922:0+3922] + a; end
12'd3923: begin if(a[3923]==1) 
	 		intermediate[4095+3923:0+3923] <= intermediate[4095+3923:0+3923] + a; end
12'd3924: begin if(a[3924]==1) 
	 		intermediate[4095+3924:0+3924] <= intermediate[4095+3924:0+3924] + a; end
12'd3925: begin if(a[3925]==1) 
	 		intermediate[4095+3925:0+3925] <= intermediate[4095+3925:0+3925] + a; end
12'd3926: begin if(a[3926]==1) 
	 		intermediate[4095+3926:0+3926] <= intermediate[4095+3926:0+3926] + a; end
12'd3927: begin if(a[3927]==1) 
	 		intermediate[4095+3927:0+3927] <= intermediate[4095+3927:0+3927] + a; end
12'd3928: begin if(a[3928]==1) 
	 		intermediate[4095+3928:0+3928] <= intermediate[4095+3928:0+3928] + a; end
12'd3929: begin if(a[3929]==1) 
	 		intermediate[4095+3929:0+3929] <= intermediate[4095+3929:0+3929] + a; end
12'd3930: begin if(a[3930]==1) 
	 		intermediate[4095+3930:0+3930] <= intermediate[4095+3930:0+3930] + a; end
12'd3931: begin if(a[3931]==1) 
	 		intermediate[4095+3931:0+3931] <= intermediate[4095+3931:0+3931] + a; end
12'd3932: begin if(a[3932]==1) 
	 		intermediate[4095+3932:0+3932] <= intermediate[4095+3932:0+3932] + a; end
12'd3933: begin if(a[3933]==1) 
	 		intermediate[4095+3933:0+3933] <= intermediate[4095+3933:0+3933] + a; end
12'd3934: begin if(a[3934]==1) 
	 		intermediate[4095+3934:0+3934] <= intermediate[4095+3934:0+3934] + a; end
12'd3935: begin if(a[3935]==1) 
	 		intermediate[4095+3935:0+3935] <= intermediate[4095+3935:0+3935] + a; end
12'd3936: begin if(a[3936]==1) 
	 		intermediate[4095+3936:0+3936] <= intermediate[4095+3936:0+3936] + a; end
12'd3937: begin if(a[3937]==1) 
	 		intermediate[4095+3937:0+3937] <= intermediate[4095+3937:0+3937] + a; end
12'd3938: begin if(a[3938]==1) 
	 		intermediate[4095+3938:0+3938] <= intermediate[4095+3938:0+3938] + a; end
12'd3939: begin if(a[3939]==1) 
	 		intermediate[4095+3939:0+3939] <= intermediate[4095+3939:0+3939] + a; end
12'd3940: begin if(a[3940]==1) 
	 		intermediate[4095+3940:0+3940] <= intermediate[4095+3940:0+3940] + a; end
12'd3941: begin if(a[3941]==1) 
	 		intermediate[4095+3941:0+3941] <= intermediate[4095+3941:0+3941] + a; end
12'd3942: begin if(a[3942]==1) 
	 		intermediate[4095+3942:0+3942] <= intermediate[4095+3942:0+3942] + a; end
12'd3943: begin if(a[3943]==1) 
	 		intermediate[4095+3943:0+3943] <= intermediate[4095+3943:0+3943] + a; end
12'd3944: begin if(a[3944]==1) 
	 		intermediate[4095+3944:0+3944] <= intermediate[4095+3944:0+3944] + a; end
12'd3945: begin if(a[3945]==1) 
	 		intermediate[4095+3945:0+3945] <= intermediate[4095+3945:0+3945] + a; end
12'd3946: begin if(a[3946]==1) 
	 		intermediate[4095+3946:0+3946] <= intermediate[4095+3946:0+3946] + a; end
12'd3947: begin if(a[3947]==1) 
	 		intermediate[4095+3947:0+3947] <= intermediate[4095+3947:0+3947] + a; end
12'd3948: begin if(a[3948]==1) 
	 		intermediate[4095+3948:0+3948] <= intermediate[4095+3948:0+3948] + a; end
12'd3949: begin if(a[3949]==1) 
	 		intermediate[4095+3949:0+3949] <= intermediate[4095+3949:0+3949] + a; end
12'd3950: begin if(a[3950]==1) 
	 		intermediate[4095+3950:0+3950] <= intermediate[4095+3950:0+3950] + a; end
12'd3951: begin if(a[3951]==1) 
	 		intermediate[4095+3951:0+3951] <= intermediate[4095+3951:0+3951] + a; end
12'd3952: begin if(a[3952]==1) 
	 		intermediate[4095+3952:0+3952] <= intermediate[4095+3952:0+3952] + a; end
12'd3953: begin if(a[3953]==1) 
	 		intermediate[4095+3953:0+3953] <= intermediate[4095+3953:0+3953] + a; end
12'd3954: begin if(a[3954]==1) 
	 		intermediate[4095+3954:0+3954] <= intermediate[4095+3954:0+3954] + a; end
12'd3955: begin if(a[3955]==1) 
	 		intermediate[4095+3955:0+3955] <= intermediate[4095+3955:0+3955] + a; end
12'd3956: begin if(a[3956]==1) 
	 		intermediate[4095+3956:0+3956] <= intermediate[4095+3956:0+3956] + a; end
12'd3957: begin if(a[3957]==1) 
	 		intermediate[4095+3957:0+3957] <= intermediate[4095+3957:0+3957] + a; end
12'd3958: begin if(a[3958]==1) 
	 		intermediate[4095+3958:0+3958] <= intermediate[4095+3958:0+3958] + a; end
12'd3959: begin if(a[3959]==1) 
	 		intermediate[4095+3959:0+3959] <= intermediate[4095+3959:0+3959] + a; end
12'd3960: begin if(a[3960]==1) 
	 		intermediate[4095+3960:0+3960] <= intermediate[4095+3960:0+3960] + a; end
12'd3961: begin if(a[3961]==1) 
	 		intermediate[4095+3961:0+3961] <= intermediate[4095+3961:0+3961] + a; end
12'd3962: begin if(a[3962]==1) 
	 		intermediate[4095+3962:0+3962] <= intermediate[4095+3962:0+3962] + a; end
12'd3963: begin if(a[3963]==1) 
	 		intermediate[4095+3963:0+3963] <= intermediate[4095+3963:0+3963] + a; end
12'd3964: begin if(a[3964]==1) 
	 		intermediate[4095+3964:0+3964] <= intermediate[4095+3964:0+3964] + a; end
12'd3965: begin if(a[3965]==1) 
	 		intermediate[4095+3965:0+3965] <= intermediate[4095+3965:0+3965] + a; end
12'd3966: begin if(a[3966]==1) 
	 		intermediate[4095+3966:0+3966] <= intermediate[4095+3966:0+3966] + a; end
12'd3967: begin if(a[3967]==1) 
	 		intermediate[4095+3967:0+3967] <= intermediate[4095+3967:0+3967] + a; end
12'd3968: begin if(a[3968]==1) 
	 		intermediate[4095+3968:0+3968] <= intermediate[4095+3968:0+3968] + a; end
12'd3969: begin if(a[3969]==1) 
	 		intermediate[4095+3969:0+3969] <= intermediate[4095+3969:0+3969] + a; end
12'd3970: begin if(a[3970]==1) 
	 		intermediate[4095+3970:0+3970] <= intermediate[4095+3970:0+3970] + a; end
12'd3971: begin if(a[3971]==1) 
	 		intermediate[4095+3971:0+3971] <= intermediate[4095+3971:0+3971] + a; end
12'd3972: begin if(a[3972]==1) 
	 		intermediate[4095+3972:0+3972] <= intermediate[4095+3972:0+3972] + a; end
12'd3973: begin if(a[3973]==1) 
	 		intermediate[4095+3973:0+3973] <= intermediate[4095+3973:0+3973] + a; end
12'd3974: begin if(a[3974]==1) 
	 		intermediate[4095+3974:0+3974] <= intermediate[4095+3974:0+3974] + a; end
12'd3975: begin if(a[3975]==1) 
	 		intermediate[4095+3975:0+3975] <= intermediate[4095+3975:0+3975] + a; end
12'd3976: begin if(a[3976]==1) 
	 		intermediate[4095+3976:0+3976] <= intermediate[4095+3976:0+3976] + a; end
12'd3977: begin if(a[3977]==1) 
	 		intermediate[4095+3977:0+3977] <= intermediate[4095+3977:0+3977] + a; end
12'd3978: begin if(a[3978]==1) 
	 		intermediate[4095+3978:0+3978] <= intermediate[4095+3978:0+3978] + a; end
12'd3979: begin if(a[3979]==1) 
	 		intermediate[4095+3979:0+3979] <= intermediate[4095+3979:0+3979] + a; end
12'd3980: begin if(a[3980]==1) 
	 		intermediate[4095+3980:0+3980] <= intermediate[4095+3980:0+3980] + a; end
12'd3981: begin if(a[3981]==1) 
	 		intermediate[4095+3981:0+3981] <= intermediate[4095+3981:0+3981] + a; end
12'd3982: begin if(a[3982]==1) 
	 		intermediate[4095+3982:0+3982] <= intermediate[4095+3982:0+3982] + a; end
12'd3983: begin if(a[3983]==1) 
	 		intermediate[4095+3983:0+3983] <= intermediate[4095+3983:0+3983] + a; end
12'd3984: begin if(a[3984]==1) 
	 		intermediate[4095+3984:0+3984] <= intermediate[4095+3984:0+3984] + a; end
12'd3985: begin if(a[3985]==1) 
	 		intermediate[4095+3985:0+3985] <= intermediate[4095+3985:0+3985] + a; end
12'd3986: begin if(a[3986]==1) 
	 		intermediate[4095+3986:0+3986] <= intermediate[4095+3986:0+3986] + a; end
12'd3987: begin if(a[3987]==1) 
	 		intermediate[4095+3987:0+3987] <= intermediate[4095+3987:0+3987] + a; end
12'd3988: begin if(a[3988]==1) 
	 		intermediate[4095+3988:0+3988] <= intermediate[4095+3988:0+3988] + a; end
12'd3989: begin if(a[3989]==1) 
	 		intermediate[4095+3989:0+3989] <= intermediate[4095+3989:0+3989] + a; end
12'd3990: begin if(a[3990]==1) 
	 		intermediate[4095+3990:0+3990] <= intermediate[4095+3990:0+3990] + a; end
12'd3991: begin if(a[3991]==1) 
	 		intermediate[4095+3991:0+3991] <= intermediate[4095+3991:0+3991] + a; end
12'd3992: begin if(a[3992]==1) 
	 		intermediate[4095+3992:0+3992] <= intermediate[4095+3992:0+3992] + a; end
12'd3993: begin if(a[3993]==1) 
	 		intermediate[4095+3993:0+3993] <= intermediate[4095+3993:0+3993] + a; end
12'd3994: begin if(a[3994]==1) 
	 		intermediate[4095+3994:0+3994] <= intermediate[4095+3994:0+3994] + a; end
12'd3995: begin if(a[3995]==1) 
	 		intermediate[4095+3995:0+3995] <= intermediate[4095+3995:0+3995] + a; end
12'd3996: begin if(a[3996]==1) 
	 		intermediate[4095+3996:0+3996] <= intermediate[4095+3996:0+3996] + a; end
12'd3997: begin if(a[3997]==1) 
	 		intermediate[4095+3997:0+3997] <= intermediate[4095+3997:0+3997] + a; end
12'd3998: begin if(a[3998]==1) 
	 		intermediate[4095+3998:0+3998] <= intermediate[4095+3998:0+3998] + a; end
12'd3999: begin if(a[3999]==1) 
	 		intermediate[4095+3999:0+3999] <= intermediate[4095+3999:0+3999] + a; end
12'd4000: begin if(a[4000]==1) 
	 		intermediate[4095+4000:0+4000] <= intermediate[4095+4000:0+4000] + a; end
12'd4001: begin if(a[4001]==1) 
	 		intermediate[4095+4001:0+4001] <= intermediate[4095+4001:0+4001] + a; end
12'd4002: begin if(a[4002]==1) 
	 		intermediate[4095+4002:0+4002] <= intermediate[4095+4002:0+4002] + a; end
12'd4003: begin if(a[4003]==1) 
	 		intermediate[4095+4003:0+4003] <= intermediate[4095+4003:0+4003] + a; end
12'd4004: begin if(a[4004]==1) 
	 		intermediate[4095+4004:0+4004] <= intermediate[4095+4004:0+4004] + a; end
12'd4005: begin if(a[4005]==1) 
	 		intermediate[4095+4005:0+4005] <= intermediate[4095+4005:0+4005] + a; end
12'd4006: begin if(a[4006]==1) 
	 		intermediate[4095+4006:0+4006] <= intermediate[4095+4006:0+4006] + a; end
12'd4007: begin if(a[4007]==1) 
	 		intermediate[4095+4007:0+4007] <= intermediate[4095+4007:0+4007] + a; end
12'd4008: begin if(a[4008]==1) 
	 		intermediate[4095+4008:0+4008] <= intermediate[4095+4008:0+4008] + a; end
12'd4009: begin if(a[4009]==1) 
	 		intermediate[4095+4009:0+4009] <= intermediate[4095+4009:0+4009] + a; end
12'd4010: begin if(a[4010]==1) 
	 		intermediate[4095+4010:0+4010] <= intermediate[4095+4010:0+4010] + a; end
12'd4011: begin if(a[4011]==1) 
	 		intermediate[4095+4011:0+4011] <= intermediate[4095+4011:0+4011] + a; end
12'd4012: begin if(a[4012]==1) 
	 		intermediate[4095+4012:0+4012] <= intermediate[4095+4012:0+4012] + a; end
12'd4013: begin if(a[4013]==1) 
	 		intermediate[4095+4013:0+4013] <= intermediate[4095+4013:0+4013] + a; end
12'd4014: begin if(a[4014]==1) 
	 		intermediate[4095+4014:0+4014] <= intermediate[4095+4014:0+4014] + a; end
12'd4015: begin if(a[4015]==1) 
	 		intermediate[4095+4015:0+4015] <= intermediate[4095+4015:0+4015] + a; end
12'd4016: begin if(a[4016]==1) 
	 		intermediate[4095+4016:0+4016] <= intermediate[4095+4016:0+4016] + a; end
12'd4017: begin if(a[4017]==1) 
	 		intermediate[4095+4017:0+4017] <= intermediate[4095+4017:0+4017] + a; end
12'd4018: begin if(a[4018]==1) 
	 		intermediate[4095+4018:0+4018] <= intermediate[4095+4018:0+4018] + a; end
12'd4019: begin if(a[4019]==1) 
	 		intermediate[4095+4019:0+4019] <= intermediate[4095+4019:0+4019] + a; end
12'd4020: begin if(a[4020]==1) 
	 		intermediate[4095+4020:0+4020] <= intermediate[4095+4020:0+4020] + a; end
12'd4021: begin if(a[4021]==1) 
	 		intermediate[4095+4021:0+4021] <= intermediate[4095+4021:0+4021] + a; end
12'd4022: begin if(a[4022]==1) 
	 		intermediate[4095+4022:0+4022] <= intermediate[4095+4022:0+4022] + a; end
12'd4023: begin if(a[4023]==1) 
	 		intermediate[4095+4023:0+4023] <= intermediate[4095+4023:0+4023] + a; end
12'd4024: begin if(a[4024]==1) 
	 		intermediate[4095+4024:0+4024] <= intermediate[4095+4024:0+4024] + a; end
12'd4025: begin if(a[4025]==1) 
	 		intermediate[4095+4025:0+4025] <= intermediate[4095+4025:0+4025] + a; end
12'd4026: begin if(a[4026]==1) 
	 		intermediate[4095+4026:0+4026] <= intermediate[4095+4026:0+4026] + a; end
12'd4027: begin if(a[4027]==1) 
	 		intermediate[4095+4027:0+4027] <= intermediate[4095+4027:0+4027] + a; end
12'd4028: begin if(a[4028]==1) 
	 		intermediate[4095+4028:0+4028] <= intermediate[4095+4028:0+4028] + a; end
12'd4029: begin if(a[4029]==1) 
	 		intermediate[4095+4029:0+4029] <= intermediate[4095+4029:0+4029] + a; end
12'd4030: begin if(a[4030]==1) 
	 		intermediate[4095+4030:0+4030] <= intermediate[4095+4030:0+4030] + a; end
12'd4031: begin if(a[4031]==1) 
	 		intermediate[4095+4031:0+4031] <= intermediate[4095+4031:0+4031] + a; end
12'd4032: begin if(a[4032]==1) 
	 		intermediate[4095+4032:0+4032] <= intermediate[4095+4032:0+4032] + a; end
12'd4033: begin if(a[4033]==1) 
	 		intermediate[4095+4033:0+4033] <= intermediate[4095+4033:0+4033] + a; end
12'd4034: begin if(a[4034]==1) 
	 		intermediate[4095+4034:0+4034] <= intermediate[4095+4034:0+4034] + a; end
12'd4035: begin if(a[4035]==1) 
	 		intermediate[4095+4035:0+4035] <= intermediate[4095+4035:0+4035] + a; end
12'd4036: begin if(a[4036]==1) 
	 		intermediate[4095+4036:0+4036] <= intermediate[4095+4036:0+4036] + a; end
12'd4037: begin if(a[4037]==1) 
	 		intermediate[4095+4037:0+4037] <= intermediate[4095+4037:0+4037] + a; end
12'd4038: begin if(a[4038]==1) 
	 		intermediate[4095+4038:0+4038] <= intermediate[4095+4038:0+4038] + a; end
12'd4039: begin if(a[4039]==1) 
	 		intermediate[4095+4039:0+4039] <= intermediate[4095+4039:0+4039] + a; end
12'd4040: begin if(a[4040]==1) 
	 		intermediate[4095+4040:0+4040] <= intermediate[4095+4040:0+4040] + a; end
12'd4041: begin if(a[4041]==1) 
	 		intermediate[4095+4041:0+4041] <= intermediate[4095+4041:0+4041] + a; end
12'd4042: begin if(a[4042]==1) 
	 		intermediate[4095+4042:0+4042] <= intermediate[4095+4042:0+4042] + a; end
12'd4043: begin if(a[4043]==1) 
	 		intermediate[4095+4043:0+4043] <= intermediate[4095+4043:0+4043] + a; end
12'd4044: begin if(a[4044]==1) 
	 		intermediate[4095+4044:0+4044] <= intermediate[4095+4044:0+4044] + a; end
12'd4045: begin if(a[4045]==1) 
	 		intermediate[4095+4045:0+4045] <= intermediate[4095+4045:0+4045] + a; end
12'd4046: begin if(a[4046]==1) 
	 		intermediate[4095+4046:0+4046] <= intermediate[4095+4046:0+4046] + a; end
12'd4047: begin if(a[4047]==1) 
	 		intermediate[4095+4047:0+4047] <= intermediate[4095+4047:0+4047] + a; end
12'd4048: begin if(a[4048]==1) 
	 		intermediate[4095+4048:0+4048] <= intermediate[4095+4048:0+4048] + a; end
12'd4049: begin if(a[4049]==1) 
	 		intermediate[4095+4049:0+4049] <= intermediate[4095+4049:0+4049] + a; end
12'd4050: begin if(a[4050]==1) 
	 		intermediate[4095+4050:0+4050] <= intermediate[4095+4050:0+4050] + a; end
12'd4051: begin if(a[4051]==1) 
	 		intermediate[4095+4051:0+4051] <= intermediate[4095+4051:0+4051] + a; end
12'd4052: begin if(a[4052]==1) 
	 		intermediate[4095+4052:0+4052] <= intermediate[4095+4052:0+4052] + a; end
12'd4053: begin if(a[4053]==1) 
	 		intermediate[4095+4053:0+4053] <= intermediate[4095+4053:0+4053] + a; end
12'd4054: begin if(a[4054]==1) 
	 		intermediate[4095+4054:0+4054] <= intermediate[4095+4054:0+4054] + a; end
12'd4055: begin if(a[4055]==1) 
	 		intermediate[4095+4055:0+4055] <= intermediate[4095+4055:0+4055] + a; end
12'd4056: begin if(a[4056]==1) 
	 		intermediate[4095+4056:0+4056] <= intermediate[4095+4056:0+4056] + a; end
12'd4057: begin if(a[4057]==1) 
	 		intermediate[4095+4057:0+4057] <= intermediate[4095+4057:0+4057] + a; end
12'd4058: begin if(a[4058]==1) 
	 		intermediate[4095+4058:0+4058] <= intermediate[4095+4058:0+4058] + a; end
12'd4059: begin if(a[4059]==1) 
	 		intermediate[4095+4059:0+4059] <= intermediate[4095+4059:0+4059] + a; end
12'd4060: begin if(a[4060]==1) 
	 		intermediate[4095+4060:0+4060] <= intermediate[4095+4060:0+4060] + a; end
12'd4061: begin if(a[4061]==1) 
	 		intermediate[4095+4061:0+4061] <= intermediate[4095+4061:0+4061] + a; end
12'd4062: begin if(a[4062]==1) 
	 		intermediate[4095+4062:0+4062] <= intermediate[4095+4062:0+4062] + a; end
12'd4063: begin if(a[4063]==1) 
	 		intermediate[4095+4063:0+4063] <= intermediate[4095+4063:0+4063] + a; end
12'd4064: begin if(a[4064]==1) 
	 		intermediate[4095+4064:0+4064] <= intermediate[4095+4064:0+4064] + a; end
12'd4065: begin if(a[4065]==1) 
	 		intermediate[4095+4065:0+4065] <= intermediate[4095+4065:0+4065] + a; end
12'd4066: begin if(a[4066]==1) 
	 		intermediate[4095+4066:0+4066] <= intermediate[4095+4066:0+4066] + a; end
12'd4067: begin if(a[4067]==1) 
	 		intermediate[4095+4067:0+4067] <= intermediate[4095+4067:0+4067] + a; end
12'd4068: begin if(a[4068]==1) 
	 		intermediate[4095+4068:0+4068] <= intermediate[4095+4068:0+4068] + a; end
12'd4069: begin if(a[4069]==1) 
	 		intermediate[4095+4069:0+4069] <= intermediate[4095+4069:0+4069] + a; end
12'd4070: begin if(a[4070]==1) 
	 		intermediate[4095+4070:0+4070] <= intermediate[4095+4070:0+4070] + a; end
12'd4071: begin if(a[4071]==1) 
	 		intermediate[4095+4071:0+4071] <= intermediate[4095+4071:0+4071] + a; end
12'd4072: begin if(a[4072]==1) 
	 		intermediate[4095+4072:0+4072] <= intermediate[4095+4072:0+4072] + a; end
12'd4073: begin if(a[4073]==1) 
	 		intermediate[4095+4073:0+4073] <= intermediate[4095+4073:0+4073] + a; end
12'd4074: begin if(a[4074]==1) 
	 		intermediate[4095+4074:0+4074] <= intermediate[4095+4074:0+4074] + a; end
12'd4075: begin if(a[4075]==1) 
	 		intermediate[4095+4075:0+4075] <= intermediate[4095+4075:0+4075] + a; end
12'd4076: begin if(a[4076]==1) 
	 		intermediate[4095+4076:0+4076] <= intermediate[4095+4076:0+4076] + a; end
12'd4077: begin if(a[4077]==1) 
	 		intermediate[4095+4077:0+4077] <= intermediate[4095+4077:0+4077] + a; end
12'd4078: begin if(a[4078]==1) 
	 		intermediate[4095+4078:0+4078] <= intermediate[4095+4078:0+4078] + a; end
12'd4079: begin if(a[4079]==1) 
	 		intermediate[4095+4079:0+4079] <= intermediate[4095+4079:0+4079] + a; end
12'd4080: begin if(a[4080]==1) 
	 		intermediate[4095+4080:0+4080] <= intermediate[4095+4080:0+4080] + a; end
12'd4081: begin if(a[4081]==1) 
	 		intermediate[4095+4081:0+4081] <= intermediate[4095+4081:0+4081] + a; end
12'd4082: begin if(a[4082]==1) 
	 		intermediate[4095+4082:0+4082] <= intermediate[4095+4082:0+4082] + a; end
12'd4083: begin if(a[4083]==1) 
	 		intermediate[4095+4083:0+4083] <= intermediate[4095+4083:0+4083] + a; end
12'd4084: begin if(a[4084]==1) 
	 		intermediate[4095+4084:0+4084] <= intermediate[4095+4084:0+4084] + a; end
12'd4085: begin if(a[4085]==1) 
	 		intermediate[4095+4085:0+4085] <= intermediate[4095+4085:0+4085] + a; end
12'd4086: begin if(a[4086]==1) 
	 		intermediate[4095+4086:0+4086] <= intermediate[4095+4086:0+4086] + a; end
12'd4087: begin if(a[4087]==1) 
	 		intermediate[4095+4087:0+4087] <= intermediate[4095+4087:0+4087] + a; end
12'd4088: begin if(a[4088]==1) 
	 		intermediate[4095+4088:0+4088] <= intermediate[4095+4088:0+4088] + a; end
12'd4089: begin if(a[4089]==1) 
	 		intermediate[4095+4089:0+4089] <= intermediate[4095+4089:0+4089] + a; end
12'd4090: begin if(a[4090]==1) 
	 		intermediate[4095+4090:0+4090] <= intermediate[4095+4090:0+4090] + a; end
12'd4091: begin if(a[4091]==1) 
	 		intermediate[4095+4091:0+4091] <= intermediate[4095+4091:0+4091] + a; end
12'd4092: begin if(a[4092]==1) 
	 		intermediate[4095+4092:0+4092] <= intermediate[4095+4092:0+4092] + a; end
12'd4093: begin if(a[4093]==1) 
	 		intermediate[4095+4093:0+4093] <= intermediate[4095+4093:0+4093] + a; end
12'd4094: begin if(a[4094]==1) 
	 		intermediate[4095+4094:0+4094] <= intermediate[4095+4094:0+4094] + a; end
12'd4095: begin if(a[4095]==1) 
	 		intermediate[4095+4095:0+4095] <= intermediate[4095+4095:0+4095] + a; end

			endcase
			if(stage==12'b111111111111) begin
				stage <= 'b0;
			end else begin
				stage <= stage+1'b0001;
			end
		end
	end

endmodule
